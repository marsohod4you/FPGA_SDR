��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�w�tܔ��R�%��«��7�:���c#�h7�u��k�u?��V/��5w��_ziCa��l��PQ'O�	C���J�#nW3����G��A?�k�gĒ��t��r5�,F�ʗ��gZ?�z�Z6isG��N=i����	x:��u�q�'��z^�m`WD����4O��E�xfG�#f=�l
�^�Q�����9J.M7/rO�?�ɷ���v�HT-�
 �W�b��Xa���a���"[�/�p�NF���_���U��j��ۀ�J���O�e �C�6T$ٸڎx�\�-O�������-�u@I):[�?��&�IE���̱'z�{:��9.W�@�	�R-�%P��X~ћ&#�W38NV�i�v�ŝŻ�O�|`�T�EMs��&fԫ�O��DK�ea��c��=g��ٸ儒��<���>�F�K�S��؍�YЁ��Τ����Z+mS�پ�6;e; VX\d��.����]aֈ��Dɕ�� jm� ^��"u�-���i#Bz�*OIs6�JE�k����r,�1��9�+_f�t�Y�q���~`h��O�evUZ�$���r{*0i�Q��X�W��R��G�W��~j��bA�ɷ�Ph�"�eetJ6���]���"�-Z���w�ŷ8�]Ӳ�Ȇ�a��w�i	�Zδ����n�	��4 �I^��vY/s�� �L���l������ԗ�ڎUVU$
���wj�{ Q�N=#��B~���w{�v<=A��e�����{�AI�����yw|��:�ɷ�Sn���ۈ�y!Wn#6�������d����	P��<�p  O��n����;�Ι@����|�'-P��R���pΛ##3�2v�er�Oם��ݍ,e��l��\���i�c��6���ӽ{y�4#O�6��)I"K�@��n��i#W����*�kb�F�=�SB}N�X���e�\��j��Ze����-�\�������]�Q�{�(Y����d�֯��V�K4�<�_��h0~8�A�2}oY�w�e"��<F}��U�_)��"+�ҥ����	ϸ#���3��,3-��:���[CL4��`8O�<Mx��h^�e�Dt|�$��Ϥ�m�+���d;�?�'��{?���P���u��
g�*��܈�kX �(S3Al�)PS�w��%t�)�e>�Isz]H˧��4Eջ'q�~��Ŏ�]��C�wh�Tg9+O�u�����u6��\
bn���x��m+t5�	[�Hv�7fϗ<��O�7���Kğ���<���!ߵUl�aŻu�c���C�����wE���gT���M �?�k&{��!���<iti�y�*I��|��� ��ӆ���;JPھp��OQ���b)���)ό�O3T���Ł,�	A�u���\f�d�J,Τ*|%/����F�Ϭqx'�������%�,2�K�k�T�w��-.=����7A�sb'\1�tg���
0�Qǂ��l��/��Kh���˅�?����!�]���ɚ�@H�-vU�a�%�:�B�`�fK�����7����>����Z�Nї$�;��j
=QqO7rOX~�����