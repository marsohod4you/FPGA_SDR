��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���y�'�>�p#�I���K��xƭ����	4u�ױ�Z�4��  �=w[�5/�)�G��t7�NN
h+��G9w��K��t	;���5k=ǨS/�ֲyb�崜����Hʜxo	YDc1¼A)�YH�e�����T���ɕ٣o�,�v�
�E��.Kf��������s(]��� oI2��Wyv��h���vބ�p�LJw�x�k��Tx���k�׎Y�_�xC����,m��������Dџ^�Y�݂�Ƒo)��9�H����m��S�P�׊�P�
��<_�C|<ދA�t��Y��C{���[���16����$�Iú:)�8M�1���$z�o?����o.W8�+J�0_O鋟$[��k&�z�m��qL��	���u��ng.�[�(᰼F�1����1�lhN��@5m�7���(�%��}�����!b�m���P:�l@�O%4����
��/�Ͻ�i�#�i,x���)�'Ǡ͜c5)Np��"�3�c���'�lg �����-�J^�������	�WŨ.���G�Q�����e�j���nS[Z��u�5)���o��+���K:���BFn��ٱ����B)�~j�*�7=^�������<A�+;�W��	%s�;Ъ���y ��?��m�;�_,�c�vU>�I��*h���MgaO�DK��0��&j��L7���Kϩ;
�]�B%�	�5�f3�N���b���5�ڡ��tN �Զ��$�n�_;���nƤ��j7#F|O���F@N �W��ٓ�>&�Z/���?~��	ƹE�t��o5Ds[�7�"�+b�~-V����V-��"��Ȕ�qM@���6d�gʄ�D�f�9�F35����h�t���$
��'�W��p"�N4����v{V��]�ޯb������ݟ����A&w��48����;\Hc�߫��O`@E(�o����g��߾�	�	8�{s&9�J��W7��2�wKL�+�Mb�jh{�8�"�qů�V��w�P���ꑩz�j!���w�q��*v�	-q[�N겔.$�B��#�M�����
�7��˥'��j�=�o,IO���s<1M�eZ�������X�pl�
Z!�Ձ�O��<@S���K�p6%w%�A�)F��n}��VU�\��r:92�X�*��U_�˩�������w��r�e���Mg����:'I`3S��)��c���R�~ȏ���.;<�,�k��y��̊/�J+tQ�e��V�Eؼ����%}C��϶��9�jPf��������tu�G���c�1���3F�{?�V�(=�E.�]��J4������}�w�&�3���$���h���N���@����4|��5 a4n��
G�����7t��U��8:����ʖ��x����ڤ���G_-�s��Ll�k���V�
�OR_7��b��B{È���T�������G�Qf��,q/�Jf�[GH�F��ZI�<!��90����'�ty�p�G�����?GИ�&xV��W�����僿�<�~��$�$�S�.RYc���Ւi�h8��GX��!*pjb�T9��TI���RؙKlb�usr���t$�Ȍ��
a~�b����r�@87��A�\B�`�t�4�tO�F�j�c����l���3�Ŋ��;zfʀMW�S'�R�I�����D�F.�R�կH/��0���.�]#�ۊ��O���+���[ʯ�I�D��VϏ�ӿ.��2�ZP�r����'�pw�=z�s9?n�0�u`X�bk{����Pm��y%�g"']���7��M������*�7\�v'�ѹ�'�]Qw��c���v:s��!q ��ʄ�ZųH
�3#�uI����X /]��� ��{ǐ�/�i�=�{���4�h??^Խ�[����ѧ��B�6dT��l2.��Vş�˱mqY|��2�U#�n�	'&NF�T�ϋ�1r˗���r�)'����,�1◠��h�H=_��w⻐����S(ɘ��|s������q��)��˅wG�Z��De;�L}�[]�ןζ^� ��94��~��G�-�U����1bo��HBy0�g���!���bx�R7+�� Y@���X{��B+�� "�����=��;T�#�8PJ�?A~����d`�����aU�3fW�ǚb|�~4�+kϻ�%(6y �t�� ���&�tKX�gXhY�%>��L�J��xǩ�[Q������<e�V����(w�8�!��8P�Jՙ�I�����S�xh�G�G`}���Ԑ��-�kA|��q*c� ��[̝I��]��z�4+�Mr%n��>�9b9�W�����0�|�:���=�[|{�Q�02�u��M=�ղÚ5�
a��`��ҩ�Ƅ�K\Q�0�^�_����\˱)-΀(L����8p�����h��^o"Ҭf@��!C�ݚh��f�ƙ�߄�$���j�%B-��v���<�M5M*�1R��0�2��<�����֯��5[%�@k�_�r�r�BΆ�8V�u���R(��+�e���YB��������� xޢ�����tg���I��O�MD7^�Y�,�M*�H|�2��}�j��'ϴ�E��Z�vRѻ����m��4z6��eu|���-]�=�F���N��Egyti�&V�P򀖰�6���HZ�ڐ�Ͷ8(v�hrG2��R-�D�à����s�����ڽX�.��� �ᡓba��J]i"){��-�J�r�"�M��7�������,�[�*F�a���;�(fdlӄ@�'� �"��ʣ{W� ���.�n>�J�q3cW��n
J�K�����Vt�Ml�D������"��	���ax�D���B�#.$��G�|I�*����"q����x����b`V9���r���@��������'b͑�w��s��e��J����[N.�l�����K!�Zw	}'�x�M��*]�ɤbH	D����R������o_�u��tCyZ���`0P��ac�lbeFFޭ^\Gp�����H����4k,ޣUs��g�l��sϥ0�2.^�~�uk��aJ��#CE�㖘G���Q?��" �F���;a����{[E�,�
EC��"'^�c�Ṹ���x�Z���׽��;�b`KBoj�#ftn����nxUp���X1�g�/��ȟܭ2��$V���v�''���p��wc��9C1�ҤMZ�%z �"m_=���L\�?^�$��~���*��w+��`�F���ΝQ�b�&�E��ϵ��MH�Wj-Ro��.�&��S<��L��"N�s<�}�u�_�!.��a��:��+�V%$�"�=��W�K�H+� .g���+�&{9�^�ٍ�F5�B����]���߫M�>�#���y�g�
�OF��l�I���@t��:e���wͫt,(DU�@����e�߮<lƭ9�؅� ��DVCqʺW��ǆ9���)s)($|��� �F6� U	�>�r��y�#5a '��v�(�=;��KB�����$]� �z��Ap����V��zb���6N� i�rA]�����lk���ls�g%���Ñ~̾�'/��2DmAX������L�bXd��#mk	�����?�k!����㔻��0U2�s&by�E#�]
=�n�	���q�yfl]���6v����V���lxW���C�3��1���b��c#��?s&���Qe⚻�=?l���J�u���$���$#����cbs;:�p�z�*�k0Nb�֠H�j�Ѧ6zP_yoΩ@��<�=�>�k�LR��}��e�J��x�T��P-$���I7V}�#��ǐ�V� nУk��;��v��le[����{4��$��+��L{-�B:X��z����ԓ��6�g�.�E[�;��*U�OD5H��K�"���T�E͙����`t-�ݭ��vsDőa�ZU����w��eYV/�Jjus�y
�ʵ.�w+7R&�̦�4�+l���jԱ^�g�'>����k�#��� ���P�,���Zl�\}����!�kA��d; �"���h r���9\<�m@�[�6|f>��Ԓ�����c��/�8���l\q��^G�:�ˏ��+��Z�\��Yya��N�����0�De�
��}u���0�V�m�i�HH��r��:"�^Tu���)��rg��]b��MĆ1�2��(���V����NE�>]�&.M���-*�0"���	�� k7$a�N(|�N`X#��+-hBVT����8?A����#{*�4=+J~?Q�{��r3�P�ȱ�K*�	ާ@��L���%所�tW9�nS�P�M�Y�������z:�#��pD/�Z��W�z��1#�� p�K�X��Me�;D���v���`m�D}��9/���OD�"j�ϙ�$�F��r8dA*;s��Qc�K�d���p�n�:�od���'&��*j�n��u"&i�"�B<G�_�Or�p���֨�����F�j�S��3�YpErV���B�,�pW�d��tJ:Ā���V����#��i��$�=�r��蔤�z�H���݈ᷘ*�<��(B��P!�w#J�����0g㬧	�H��o�z�䖘:]��h������H�T�p�� ��oM�r�$|�Ѭ���9�R��꘲��$�D��ř����-T�h1��GR�WE����JZFI\D�Ir����fL��99��yNz���:ҍ@�6 ���G�y.���H�9��']��<��{�ܔM������I�P����G��-�|�OJ��|컵����׹,�iYQ?'����86g�g���`(Yaq�8��8���61�l.����3�cM��'��;�ݩ�*��L�#�wq����;@�+w�������e������k�	a��c@u73\��e��D������L�:2df���W��,�8�� �j��a	��)�[�}P�NG+}N�f�#�S|9�)�X/Ҍ
�"����n0�C��tɪ���S� ��#�xjޞ���	ܬ���*���Х��tr�l�ʚ����1$�`z�N�=���l-;@�5��`�(%E���P�5��[�<�e�O��n��ږ%�d5^�x�2��㹝��M0�]�L�5d���D�}Ly[ٰk�&��$�mV���N�ytP��.L@B��u�ן�6s��X	��uf��t�z��5pAP'�>,�A2DL��.|%�$$�bٟK�4<�,4������PGЊ5�|��a��(Z�>Y�M����W�s����$�����a��zg�FN��0����r��i�LX¥�Y]�e��a��@F3��`��EP�'�P^¦9��x�Y��]�B�[��K?2�#h�{9 �^��{�1³�6���cG]�m=F�e��ڝ�cea��I!e��$�2�/�ʐ�F��7Hw��%���սn2פ:�b����m�q��2o�C=�M���67n��
2���r��'��J�:yjR��(8��M�+uX�G�Ufk�4�D<�5��RhB��f�Jہe㙙�C���c@8�)tᗧ�f�T��>��A7����tX����2���^����ڵ������'�x�>�%��5*]����q+@6�֕���|^m�D�����%����� �t�L�����Y�g7÷6��BB�� 5�o1y�@�|�rE��a��!� F;.�HѰ�5ɩ& œK
5������1����bf��:�)���PSqK{+L���k�����R�<F����HK`]qpɆ�
�^4�u���(ya11Ò��J��sS'�BmK�
�eE��b���1د�H����%U�����b�3��4'tO|�=��*����Y<�<}�.n�έ��RN�������}���|��U�H{1�N�&!�sB��h�Qj#ū��Z$N�	'G��[uF�|��Mܹ)nd�X �vҗ�T��k�D��Au%QN�p�b
�=��	9���Ul|'���uqc�>���7EH#�m����a��&UƲ߰� ��0����}U�Ώ������pO��q����}�My���I}f���]�����n�'.�m��)Z욷�#�t��E_W�7�
�?xn%��T�F2Kj����A+��:go�xӄ�{��4�Y�`w� �sp��R(,UL.���z;ٴ�*NN&@(ʪ5�U���YP·>��Fl�$؏������P~�J:�g�ST������$'I�vj)�E�g��wdCz'���]�UD�UX� �D������@t� ���bH�E��ļaS������̖a�d+UQ"�mT`b�,�^��jy*
�������qJ�AE���zb�����*��~U��&�4��D��h�Cw�� �Z��z����|Dnm�Pۇu���>�1�n!�~Dyј���n��<7N����>>�Q��L���5i����F���p�ɢsrqDV`A�-R��V��UR��h�m9V����Q;��E$Ɨ$)����u�q����b"H��3����n�&��w<XZ[�=$�k���>>g;=C������D�aYggg�G��b�L-��5R?o%2s�P�&vdP#��h�}��x{i$nl���k��fY��Dþ�";	��s}a[�tg�����*�-@�k���
p�w�H��j�㱈��BC�4�Ǵ��+u9�W���ĦD,����3�
��s c���.}����)�FAWX$+��t�{��h<h�g�I;��R.�2Jb4�KCN��:�J�X�H�1��?�	����y�q����LW���bc��hҏ����d��6i���(�1�VM\�HI��@rW��z�rR��ts����gx'UKH�^+�˶5��'(�|S�� #WKs�>��^P�dg�O�g�}m��ƴ��?�4dm��9�����D�1�)q�7ր>'���˧�Y�WU��m�;��	6������.)�~�(���ciG<nJ�ku������g�+�@��ܮ�s8��_kf�0	�K���7�=U
*0y��$;�������J�/t�?�٢��J���<��w�_��4�p��!Tcvϝ2�E=o�s)\d�pb͍��Lg�����$ᒾV�KȸR�$Zz��ۼ
�O��\������U���G���U�n�Q,,62 }4��y}�%�<Q���P���Z`&/$ i/M��k�tfu�L�Z��
r�'$�A�0��D?����w�0��{�{�:M-���0��p��<YL�,��#E���:�a�q	zI�ٖ�ɦ6P���r��J���%�c"'4zKΛ:[1�
�)s���՘4���a#�m����%G#���ME�ܳ�#����%!���9om:�j�{Uu��A����TH�lBR���0�������ű�|�V�#�h-h��$r[�P�?2^]O��گ��l��jz�w���t"ta�3Q~����z�94u�����gR�̜=xX���!Fσ�wh��6%o>�ŵG�:}�%��{�U4ӏ�����i]��k�RKWm�?4��M�쑁A鴱���]�xts��$[���*2��!K����T��'�~���"RN��z?̟��I�S@��Τ����r��!�D�Qݙ~cJS�7�M��\�/�ԇ�h�i�� Uvb�~��q�o�U���|�vV��K��a,|�'@c�)tN�.n;z�ܡd��S�yxy����(ع����0B/ L�����]��&��7�N(����uC$䘳�NS;6���ޢ㎧� S�����n~d�����%������$�$���;�Q�'�D�8���l�~�����:�(cJ��	w6 K؍c�y��aF��X���Ő(� �F0+�w��h��0[$�h�`	�I����xy:������e�a�s��]��*į��~yPg{�D�\�<���:Cw�jO?	�!B*./P�(�l�o< IǓ{�.��B��(њSj�$U�}��G>/��(��/���.��σ�ׯ�'���>��v��q��I=)���"RTP�j�k�nꏕR�����˵<Ʊ@���+��`1�mݙ��l��]��	��>��&��C�0F"�%8*.�T��;�LS�q��|Nq"��
�	�.�SοV�6�Α�^���eC��m\��Z#j�7���F&��+���;=�&������l�j݋��=Y�K ������b�%�ʢGig���&��u�nېn�w��u�����vs5���F"�m����
=��t(��A� x��H�EDz�ߘO[̍}��냠�e���$nS�(�
ТY߾�Y_���:<6��w�DZ�>8�&��p�4�k���xmm�ߦuӐ��im�a���:@�������"���
��ߣ:l�=�#KY��h�ߪ���&�uZ�Uo���S
.�
�Hcu����� ��?����)SR�����o3��B8�҇�<P���%�?x�a=�+hb�D����Ȅj�^j����=L_Zw���TY�w�C�N�H6�U�u�{���Q�"�_��V&�Z�v��o�쇏�O��a��P'v����wޛoošg����O1�l)b�L|��F-l6H�<t=%���>D�r��
���:88�;E�{���
���<�vѤ�ѥ��R��f$���O������Hcw��V����������O�zE���!S7A�h�����������zqI�X΍�4��*a��u� 
�8飗Z��1Lrz��C�|���� �`9w���	��ܜN��T�I��5��)�T���@�\[�+Qh-��	h'�홚h����QC6�eO�͵AZ��?-��2���^ʨ�!�����j��YA���E�n<�!)�v��Ԩ�l������.�s�$��6iq�|G��8��]G�;��ݕ�EXq����U�V�0zt��6x���߅�ˇ��O�dH"����;�7���JA"ӏN蟛�l�	�{ �+�f<4A}q��S�-�n2O�����{�#��� n#eF@
~F���~���0?jX��(Li����bc;^'x�އ_��D���W�QN8�D=�������^� w1t?e��l	�8�yw���\	�aX��*K���&���	���w�\���gڞ4��l���l4���,�����pQk,�5DB|-�U=N��آ7��/vi����f�F ���n)��)(>�]e2��T��>���Gl�Q��^��=a��x����D���&����?&���6�ޤʂ��X��b���F}f�^X�A ��$`x�B���m/�Ao��tχ�)FH�J�i��҄�e��Z�C�TR$�����t/�[��^g�M�^����k��j]Q�gIYK��-�:y��؅GS!����*�`�jd��F���30���2���2�d,}h�/n�Y�	���V�],��S������Jt�;{��k��ɝ"�<8f���]� �L�O������ǅ�������TO;an�	/C�D}���Q�Ճ�'���񐠥��뮱z 3���5�RhA`Ǵ���r�3k�?�$|�l�is��B&��=�/����S���hf�׭
;0��vE�y�.��}��\�z���� '����Z�<�Eۥß�B��s<\�CH�J/���u%�;6�\�?3��4��{�WO���a�{��B(�����)7�|�
�]�N�J�;�И�@�ʰW�	��3�pV��a�s�t�I����]\,$_��'P��Z�g�#Ofv2�N	 +m��׮�^2׿j��"��ξ���� t1��;���� ^�q�N��-�OB���H��:'���=7�'��_F���V]�{���el�Ɓ(�i�SW��&&/�����B8?�����>�d����]���t�o�ϻF�\���b6K�,�>}��୪�ʈ���7l���R�:��|�L�mcl�'��K0��.�m�u�v#t'$�ˉo���VD�N�K�kf*������ A�;8��O�ClRn č����`��{]|g/t�x
��l�ޭ.�eF���)��d8u�Ѣ"�cm���2�e��(a�V%�Zbk 	�����Y ���CklE�Sa�$�aGV&�I�RW���5��/a4��uݳ���ݛ�.a���f�6�jRM+oy=2��`Z.Ҩ��/S��	��#�|��$�[��=�9�8:�4�9�;Lv�}�<�����/����=�Sr6yШ�ۚhv�F����ҿ3F-#읋5�<��7rƔR��2��J� ��<DLI�^���f�r1ǎ�!g/�y���ZA�\�U�\�uB��[��J���44��6�N{��s��� ���)+zK�`'{���Ȱdm�u����'\7��40I���.���L X;�8(舌���'����A�\��]<JJ՛]��Q�/#)����,|h��8���������&�y�LJ[Y������X ^-$��p��ԉ�[�5ooɌFk"5��w��:��|�2f���6ҕM}1di6E�7�lbv&��t�ǣ��\%�f�b�9��j��m.�zK��L8`��d>�h�lDf�F����)�wN�����Z�Km%#EZ{��y��7/x>�H�p����0m���w/������[!�td��ﰞ߼�������Ra���װB�m�h�>6��Uɔi�������n�;u���qz��X�86a�%J�`0������Q��<�66�?W�v�ޏ��Ƭ�↱ό�rp�v.dW��"��V��DP�b�}0Bl1�o�3P��{]�d������F�m	��ޓV�4U�e���8�mjv����R�h3.���>���� ;x�4_?$X}R\�EK�Ǜ''jjC2���1��}dH+C�_�����~ EQK�>2�mSdӪL��.�a�H���ud��t.qY��wu��� i>�j����H�}��������{`ʆ�������ʣ��aA�g���Ǫ9OV��[�C<̒�$U�ll�΀�5`L(>�=�p)1��<eQ._[^���%9����E�
���������3:��f9�����.������a5���J蔻�l�2�:�D��������k F�{�+��������VfU|��gc&F3$��e��j�VJ>�� %�|[���^"����7�3���a�*��;����5g*g�J��꾚���|i���-�qg���y����I������-�):���@w��<]�R��v���Ae:36�*PVVR�ﾹd3��/�&\�I#]{�J{7#ߤ(��<(1���R��p�T�α���3�c�H�ϟҿP��&�� ݿj]x�M�����L_�L� 3T3iV�2�Z-Y�Y�{1/����㭛)���}�VU�?$y�3?����e:(��mjR7�F��G=�W��Z�'�N'�coÊ�
�m��y3|6�-��d��r��Z�.6>�S��PB>c�I���Ү�;���¬�F& �셀"��-��Қq���J�EapE!�鋧Y�@���Ŷ�Ң��<?��0��ܫ�t!�Y4a//;C�����H�i��YT���N�q�"��6�Jx�w_�ct���E�/�r���:+��n+�� # �o���Y����d�U�"�>qB���8��(ŧ(�se�R��AĴC'�#��! 3�1��ά�O��9�e�O6�s�
C?}G�Y[SW�P��r5Ѹ��Xq�V] Խ���Z�A\E��)/�!/�,�ļW�9�?�vmД1�-��d	N�OI�7 �b.ѣ
?\��	�T�%��d�qd1��h�ظY�C&e~��)�\��k�)o��\���YÂq�#$V��T�젓�T�R�kEP����_�j��e��2�}��V��]i�ޘ&H�		�H�D.�6y�Jd�Ibol���?m�߀V8��[�h Qȯ�Ʌ�N�r�B�v���ڌ>BÓ�,T�`W��33�*�y�]��Ո5���ц1���~�/���#��2�~%x�ܡ����y��� C7�YvU����G����Ʊ�P�NEs�1�N�_a��}8?�JM_�/f7�Wg|�{�Ϛ��������O�oIvgC�Ջ�?f���
�*XG,�t�`r�?����=
�]H�,��q⸼]��+r��37�5�����R+�1}j�D~P�FP�.�q!!l}Ϥ�� @�(��26������xD�S�z�����|\M���� �)h�k���.ɦ��{ �K2B�o���z߶��B<��M'�̕�ҵH�f�@s��n~h��"M*����J0�2��;�g��� ��]�_�*<�d��!f\k�z�YKϻ���f��Z�Q�pX)d��6�_�4�᮪'q!,��
o�){J/p'���O�ZC{\�d�w��H-� ��.р������k���em�[(�<M�.}0W�I'���n�[C�9f�x�0�A:Z>�����?cėB��Z��!s�s��
���'2��p�
/h��6JMyZ��c�y'[��7�K�0�Jd1��WY��ʍ���� �N�?��׏���M1縮�������=��{z��|}?�QKY�R7����7{O�� ��@��e/�UH�a�����fK��dA6��P���6<�t��� *��I�H���B�l�_�gW�MZ^܌`G��F�T4��n	�d��le!������l���IRh���^�9�]?D��G��ʹ��)��ctW��-���3��WmC�x�(�8�R����jh��ė��􂄱┰{�W�Id��'pW����F�\%���՝)wy���W�pz�mX^Y�u?���ڰ��ק����k���\��4	C���<��o�+���Q�̥�εCm��*�e�X�$-�!���)�A��i[�����c�X����m�%8� ա���� M2�|%��WH�.Vj�\9W���%**��� VV��]�����i]�o�}��,h�1h=��h��8�m�:א�ڶG�������/0f�1~М0�ZOc�m�l��|��D�D����R�5n�K�߿���L��ZC��{�Ƣ�(��	W�0�+��G��FL�"SS��~߀v	��b��߸�9�S_��ő�c���vq���:<I�d^�h�;�7;��c��]�����F;��ʲ�;�������nh�~&*qN�w���{��۩0�1
�~������3ă#%��)�0/�CgZ��i �'q��0/j���o�l�J$G¶�KH)JXbty��2c���� �Ld;�F�b�s�]�D�X���\P!Z*yI��f�0f0�MA�\Ǵ����ږ�xRv����:ûȖv�h��Ո�5��k�Cy�2^���mϚsge��ҶC@(?!�ܗ�@* ������0�B�7��6[`O+�b�j�"�8�ݬ�B�����%�-2�8��uda�V�����|,}a�+U\}�A�\Ӎf�IKz�so �<ȫ�O ��z|P&�7��-G&���~�<
`p�5���uy��Z,�9�z�!��'?��NXe��<a{&��j�%F'�+��*��џ�&�?�mi�B;�)�K��8�T���Ў ���[	�+�~��B��)e�N�K�E���s����wd�S��C�H>�Uc��:x�@������w��՗ZY�*M墴YKӜO�?Ä�T�8��{I�?�6�Q�����02�8æh��q�l��.�)�+|>�K��{4t�ܻ�_s�Q��.�"+��� �-�>���I(�)�0��8�)
����m�P�Y�z��L_�R�$�O�����6^�V����ĩ�(rf͈M��ɃY)�:)�s6Av�|��ڎ��N�g�6�V�t���,�o����.Z1.
a3�ή���G�Q�(�L!��3�E�[��qO�� �X)A��S���8vv�1rn���O��|xdE=<�tx�ҙU�����"�	��۾�
PW���O�7ָ���[�����'�/�6�4��A �7�^���T)%o��F�kF	1�̮��n�`��~P�h�^1Ĵ��H�y:P��d�� /���VK#�$65�)4ȩ(�P�eW�	�Q|���ϑe;����`�6QG�K�rN�ڄ���ֹ�N"_\3��W��i(��������%n2޿T�3i�X2y\��n�*wп�M�=�$�3����-	C%�룊ܳw�~l�B��g�������~(k�=pC>L6��Y�s)����6hio�yy=jl�/ˣD���ħFw�D�g�cWZ�H5/�>�>��H*A��U��*��|N@?�U�Ĺ���,���7��7������8����!� �%�?�"��-��O������nD��w�r�ے��B~�f�;	Ƅ���;V�(�Z����3��OW���'��/���P惭��L<�F�6��Z����o1�w}��fO_�E�7�ރ���D��9bXL����l�Y�
�8�˅���+�6��c�T# �ӭ����{/�p'�-���[՛/�C3��n2�����bԂ��!V(]��ǊtU({խ<#�O�W�y}Аf6�W��ֺH�a���3��U�Pr�|
y�N(E
g�K�v(I�
�q��L>��4׊�:Xp�*:�u�Ԥ�J3��֛��\����b����\je������ɢ��v�6R��(U�ID����������W�GEx�ѥ�����#w�+8kb�^���آ��K~�R���U#��tX7�	��`��X�*�K�6�������o����`:Q�}O��Z�?&��'�D�#��0��2��t�&
N�a�B�����k�l�-+I�����p����Bs��_w;�nB}oI���ns��5K�A�Ew9��/�_jp���=Mvӊa3|m-��C�&U�E�C�o��	��)X2{F��j�|���G3�t8�a�,�9y�.�����<p�]c>�l/5�y͙�[��^}(K�ܠ	j5����i5��J����ι��?=�K�8�)�+��
ಶ�@Ba�˭�|<����_V��!�_���"�2��+�� )Ų/������t;3��c��d����x���ҐH'7��
ǭx1��f�E�6�d�$�lq=�� ;�"�96�H�>p�τ�菆}9��Z\��k$�{�����Y`��>�	�\�;�0$FWT�r��՗�K=_$�F����@H4k��x�T�Qa�J�5T6����V��S��𘾀r_74Y�v���j����,���;���d���dVs�X��Q��$�T]��4i+�Q?kp=VDa˽_��aMs�n���"�k�����scƭ���Afũ�n�i21tR��%�'�t-,��~G����,@C�%�����$��eW���m��Z����X�]�b�=]}�!��l�홣v�WBs��SP�Naƪ����i��̻��Ș��������.��&|�Ú�W`�^O�����/@O���|)q���#M�	i�-�4����:��ܞI�Y����k�s����L�u����?�o��^�ΕGȞƤ�;����Җ�X���"�v�dC%:�':C��}[�cl���p�#87���1Hӏ5?��#N�axy����,r�:��ա
�&YLٵ�$O'��1مUG�P,���T=A#�K�h��~��<C� m��a�����b�W{`��٥_a4�biff>�9��(|p�Y�Q��6�6`ÕԞ�,$�W'�֝
&y?m�Fs7�K{_L���g^4�olmOӼ�������f��J������HH��伥��81o�%��[N	I��M���wv�#}�S�3 r¨zZ��6�X�Wv*� -'<� \�rC�F�K�gX��n����s�s��!���@c���h�	
5�^�p\;8}���4/�I@���P����U"�l�s(fg!�/	 d�Yf�t�<�"4���*�UwZ԰�_<�&)1G�qD�H�K����p�s���������>�WZ]��2� ���N'�fNɯ�!�VE�15c*�*;ܿ��ٴ�a�>�;�E����D��������[?rr������Ov�%NM���e��]���x����Lx|4�D�u�;��?���iӈ��1�qx@;��Y��.�x�M��;Ƣ�<+�0��Y����:x?�˨���!��+�mx��/qx.��FRdU5@Cr�Pt�]w��c�*�D����8� k�}�l4#b�)���$v��wn��]��}7���4eol_J���^���_��Ks�����˱���"�d c8z��t�u9V��L(O�o�\~8���<������hs������%��S8���̋8�Z�<#�wk����?��y#`7ܑ��ۿM��~��<���A � %j^�I'ai�*�m��-�����=�^M�ހ�_j��d�ϸ�y����z�׆˲8�:8�wRN�-?��C��R�$1E��qb[y�l��L�-*��b���|�5�H�v��g����R_$�B, ��޴l��Q���8�3hl�Zϥz�+����t�/\�.�zo����Q��5��:��#�%;p��$��ك� �(�̘����� ���H�N�N�}���A�֎�d�Ig��J�27�IMqfB�h��Ͱ�9Q��2���j��������ī���M��
�'�`1c.ĕ�N�	���9?�wf�9K
u�[�d5���o"X��*�V����ʚ����M�'u�2���ݛUf�St�a^r*Nҡ�/85�׌�K�J�?_�L�Y�[��q翖o��x{���}�z�ͳ��5��4BEQv�әq��cd��)�t�('hcǐ�klA�ػ���&F���z�G�Da蹊D�ڿx��lޣ