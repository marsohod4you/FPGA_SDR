��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`O�u�_|UZ������CC��T#���/[�R'��wZ���4�H{E<K��ۡ�?���i�!��,�bwݍ��]C�t��b������ �	a��@�"J(��n%��W�"��=C�,���L��%��[�N�[����
aifA-����?G�b���:��(���\�Хp�l�+䒀��d�G����Ѻ��4m ��O�H+�S��  ���a��i�����طaV�%K��i��|�n��d�l��k9`'��+�ѡDQ4�`2��n��Q�*j�T�#��x �o�t)�S�O��UQŏ�!E���m�݋�"��$Nǁ� ��>�_�x7�yx��6!<뵧��~+ά�X´V����Ѯ�.S���e6��L�N�������[�"T�R��^;/;	�y�뉩�cp��'�;�T��$�U:'�Wk�S���[V���Xx�aT[k��P��we�#��,ׁw�v�q��#Pׇ�ì��}E��hW�i?�}��7L/}���K(xӎ��(��Z��q@�J�&��t���}�,��e[w�*s��6��4��/"ub}%��E�"t����I��.��@`I�a"���W1�'R�q�`2�����u��U`��_c����i�_g���I��k0��������7�� 4��2���n��&o�X�r懨L�a�2/���.
����-�B�/J�K<L~�2%ׅI�9�4��"0�$��t��~�m@[<��¬b�AF�\.-�}�\d�|�o�	t$u|�_5�7nV2���1z$"~ ���*?d6����ٌ.b���l��
_	ʇl��5݇�s_'�j�("=o-ja�r�N���#(�&����U��frs��u[��g������j���O�Ҡ)O}+��� �7��9���t�Uy4y��5���D>�㋺/�I�����d�x�'(�~/�wE�R?$� ۄ����J��#ƶ�1�7�s�3��5*�>���~U�1�⡘��Sp�3�꯺�3�� �vSe��b3A�̕E�>��}te�!GۥP�J��g�sʠ�9�.��}%� ˴t����=
pd pW-+A�vm�	�����Tt~������F9'9�����7��} iXWb���?&8_� �2P�GN����Wy��W@�3:�&㊰��%��c��]-3.�߾�!��k�/5?lo$�� �H@#��L����%���>�G"��rqu��::�83�ä8VYqta��ݪA<�u~)xH^�hO,x��*D�ZCB��`�V\P�ȭ�u c	2��Ns�ǘ���J]�0{5�a�~�5�#^mt��*T�s E$SE)#R�AF��D��jw䌾��&&�A�Sn\c�s������f�ۦ�-w�Zhd��a�/��=#�J�ж9�?�YP����+���� �:���)A�yRu�\�3-��4
j"��Z�'X��F�&���؅���X��0�}�)�>������;�<YMW��40=B��g���m��S�H��hG�U�]۶���Qz�����~�1�
�h�@<�q O؍ͫ���@��d�c�W�-M[��m|隦�����UI{T��?�܊;�9�������Ծ��Kkȿ�����&�܂��Q��Y��M�+�?P ���4Ai`K��-�L���04���m�r<�'���q�^o��#(������6 qG����aA�9�[�hv�v��[{`.ET�Ό��3���Z��OI,��gă�{�WFȊ�򭶿�A5�F��<k�z��R�6���+�/�SQ��,�2i�E��dwn/�)pX�J�Ǉ��$��{2��C,�	�֘,e/��ՏN^�#��̴��Q��7�*�|�Y���`G·����:w@3�S��Z� �5肞��Đ�[����Z�J�T���`����[���'0:�	`�d���8u�6�oFDV��^ӻ�P4+��)@��X����F�����آ��|��S�ɦZ� P
W�-�k���J��>%�i���%R�$�f&֤f���J��_��Z�\i[�$*^�v�X���Ӡfq�#�\�u����9�	$�F�4u����&�>~���������U�z��Je�E
O��lJ]m'JA��ߔ2�R��,�ªМLU�h�z�����KB�aeb׳�1�;��g,K<�!���K��ە��zk-q���
#��1�ζ(W=7�.���0�@g�`�.x�$$�� ��YhE�߃yq@4nl�T49Z���\�U�1Q����D��Sh�`���������Q�����d+�Wdڒ���X��p�h�f#mOf`���ng��U��s��+���tL��Ȍ����I�0��9�	�1�#�;[l������- �&��;��Ë�I#>Ե�9.�c?�4���v�Ալ��I����Mp`�)�
.M���Z'xZccvV��H�3��,v �@R缧o�"����q~R�9�pM`��,��8?ý�]�<��1NQ��_~�2������M�h���s�$� �w�9��:����OBL���}Q�%���C��p����f��g�1X7�{��x��G�i�*����T��_,�R���]���U�'��J�˫�+nP�ꥪ]zP��@�ކzT2K�)g� c5U��G�gl
Z�&�9���G$���w���ОN[L�q�E�`40"�y����J�ҭD�p�ꈿn䘘�&��8�}0~e;�V�}�/��3M��=�$z3���j���L6ZGb�-ad�*Z�7=�����j�YG,�
��Bz٭>��,��ۺ��M����v�^�F`'�[�1l�.t�PK����KZ���[E�~�We"5n���6aRVuܫ��Y�&���"���^�.�����i^F��W@8��HW�fF���r62+t���(�!�\Ը��wI:@6�h���C�/�� ����Ft��%|׆��ڔDС�:(������ܩZ[���'��9��:.Y�37R���b�q�$����Nfؘ����ʭ#)W<�� e�(i���v�٪z�z)��|��=���>*s�=ۡ�[%R�:����R�T���/.�V �=H ɋ+��4��F([n����!/:��"5�Ӊ�;��J��\��d�)�o۬��B������P��$@��y����%���,�;A��k��f^@mih�rω������g���>�r%b��]�-8�c�=Ñ�̻E��?�����,*�#E�:h�2V�����-�s2�Τ�{)'�4m�|N ���Ѻ�@��I@V��#Yg�-U�2&B���gX;��#�����qS�le����@�M�M=���QDP'+��51��{x��n���LF�n��w�{�$������oK� '�;���Dm41]����1&̪ͅ:~�jqsHl���u@��B��j��c���{/@#�R)����u��^M��xS��.�3f`dU����Ñ$��ծ��)���M��r�����s�̼l��>�PX�P,�/0z0�)T�����hM����{<U��Zʒ
�~�-�G@�v'�u��ͭ/-�A"�:�p��d.��j��t�|�x6��W/��(X�LwYpG���v�Ө \y��U���-O,�$��K-E>j�/2�6��r�޻+�B��HC���t]ۤ�Ѽ`��!��-�B�MG\�wt!(dP+(!�#��%I\���ɥ7�&]aP�E��h$n�reo"����a��)��G�|�Yt
�ŨP�d2�"�J�<pܺJ}WS�;�ŗ��݂�P����F��G�ۛ��!�~&9#b\�8\U����L_�n!�N����q`]�b#�4��8�}��1j
zu��Q�jN۵$�O^"��1�rX]�Ĥ��2�?����z��Q��Ad�'���UF����6� q��X��'�Ɗ7xӞ�$��7F��7��7Հ4�8��eȄs�Q�v\��eҒtB^��=�p+V�&i|�!j��&9)���	�<���qj���Z�h�����^�G�
-a*�g���$�O�῜t���k��1:��W�ȷ8K��hiq~��ş\���Ё��N�c5_V��S@㠻+�G��+��^M]f0n
����E4���
��B��M�\}+����:�1�v�i}?8��6sl�
hd�2�m�fu���P�Z���E�9.+ö�-�=�_BOm��y F\'0�$� ����ȃ�V�]�`��|��Δg`դ������2�k���*:j;NJZR�c	z��\���ji�mh��b^�g}/�z�C�.�dF!0'Ƽݗ�JTWKի�h5d�o90�A��/�_Y�i��(=?���*��j�t��x����"��� I���b�KZ�ٰ�>{\t��	���W����Ur����kI���o^��͊�����4N'!O3�i�y>h����Ҍ��EӠ~�,���M���R���N��)�ȶ��TAd���U�&�ّ����F���؏q �:	ԏ�D�d�Cу�u� ��Y��>$�����~��I���i�0I�d�������y�f:wɶ�
�F���<DgС[��S���o�S���ė�X�t���B<j�A�V�^�_��8Q5.�ᛠb���C�<�D�a�B/̌Rω��xq�3�0���-��L9�4/RB�p2����e��j�I���I��F`�+B�Y~�!���(ة��
��iD�J�Afx��%b爐٠O�&�x_��K��j���ǰ����*G�wAY�#������m#���Ynh�j�� �0�N}�Qs�����RWE���q&\VZ[S4���T(;!]�� �L�+lL�Rd|���*�S����]箅���>�����RD���{�d���O�0}ۇ� ,ʼ7�q���j�ҕ�m�ЦV"�"e�>D�y�u?�jEQ� �$	Q �ݱ/��MA9L,�߇w⊴�螂� {�n+~�(ۊ��=HG��Z,�7��y�ޣ����q��C�1�I0jOI3oD�|,Q�Pl�m/=�����D�=.`����D��� �C�*�\ִ���q��tmV%&��fY��� �$�nJ��ܸ��<N�8���'`A�P��Z�:R�@�9Y=�I�.�W��O��V�SQų��5)`���u�M	5_�V�=�Of���"3Q��T䨆#�uхr����ʃQ�j�+P�ӯNӕ��sճ�M�J��F�C�ӏ���*�LO�@��3�`_!�u�l-b
;��E6-�/Pa���#�S��$��%E9:�xB�Qϐx�v��`�,"��ل9�ooJ0+�&ވ��ﲛ(W�@��(�X�����!<��j��o�:*�� 2F]��pf�%�r1��S�-D�;:�l�����p���{�����Z��t�4x]g��z9F|�K̪M�wr�z
`����W@�Z�g8;p�^#$�?����X�q��D�_&�,�<���-����9�����nf��UѸ�{Rg������2��I`�D 5�nh���$�?���+1�P��gU p��)��3� ��D���)���Y�P��*S�a.ٺ�h5�V%r�dJ��θ�Ū�Hw�M���|.s��˴��[5l�t��]�H���P6'Fe����S;@�KW��+���X�W��k�4"��%[�Au�T雾/���	�b;\?>��E[	��g�Ɍ�X~,���\��4�͚�uw�
M ]�'��חe�i�솃��r���ۮD�  -�?�yP�G�gg e �TL�&gH5e+�ã�(㫷�{����炦���)�ݩ>�F�_'�L JգfYtDU�&W��"#j��Z@- r9fU�堢�tPJH�0�'�-��Q���|�"���XЗd��@����ャ��bW�F��V%�k��i�����`j��~��_J];�F9�uܛs�/Y�|�ژ���;��:[_��f�VH=��Q�'a�LCX�F��|K���EY\��R
�a~�1O"�p�H�`���G��0�o�ҩ ���:�r���d9�����xƾ;2�8�X��x�k��&'�#RS����c���R��A|�z���_� ]�-��ֿpn���5���+I�=�M���RrR���������1������\^IavO�0}=���M0���K֑���!9�ըhD��������?�1x#����tq�.�C��ۧ�b����g,}��FN��*�qS���pѿ��*���4�8�de��6m���d�X�4�DDK@&�9?�����!d�%�av������d���.�_w�UHD۶��N���(��� ��ɷ�C</}8���{���K���FZ�\����̡��9é�+�-�Z=Gj(��!)��ޣ�� ���S��}֝�5�L���́��oP�/�!�Nm�o1�r���^,�C+���jmMH����.�zyF ]���6RD�<������U1[='/�z�M�dX��k��V*8�OTA߀K�z���9��'3��A���3b"SW^^+�}��f���w�\l�؇t&%)��b����:5��0&�i�K�7,}��Q���a��>���C�f +�[����jZ��skߍlK�s5I�;^G�x�GC1��3��b��	m������
_ �����o�Kl�j�R���'�wXv����W�и0ˤF ��� F���:�9^uNb��&֘u�27����C'�V������Qي�B&�{)}�e%�ӻV�ʺ�P�C����1�L����>e"����O��WA����Д�C���`\{�� 7����d�ꀻN��?���6g���g�A״3�8���O�q�y$����:��
����濅"���ó�0$�cjQ\�49!�Ζl��ҫU'�~tX�.v�+�la���r� a?p]�=�m]ue]�>/�`�8���E
���F:ل�d����(6��E�F��E�����u��N�lDMJ��q����ޖ^�C\���c���b2���7�ChaX�KjU���Y�_���R%�×1���������P/���zd�s�E�Z��=�Ӱ=�� �9�{,9�͂�ETKaj1nOz�iɍ�B��/�S/ѣ:�zҘW����	8�8��ѕ������
��k��f��^�)��ɝXOJO��p%�{�Xjx9����n-Y
}�t�.�-O�6��q��bm6V�<Yv(S�듦2�i�Y���&��)�z�F�����Q@��9���(��1]�_�5R�P�m�T	)2]�5� r#���!�cjk"��+��jV�g+D�e�笞E�����G�э����*��+���u����}�[D�}�{ES��V�D�~uOH�j*_�Q���yf��[�L��gp�j��{ӣ��U�#���A6���xL7u���z��j�@T&�)���(gyQ\����oCoG���`��1����H#�[�D&���'&c��X	z=z+�(��@[��S*��F�Va1d�! ����n��8x,I)�(�N(��|�)�Y7T��6@���Ȕ����P�|5�Uk�⡂��{x�=�r��}����W>���'Wj۞G܍���"ߨ�W5[�����{Ӹ�g<V`Q|[�+~�.R�5���d]�W��x��R2�L�Q0�V=Uc����[4����zS�I���/��ޕW�ȳ����i/ѭ���wPxoš�e[�
��QO�]p9rƯ1���HB��R�NV}�����(�����Z3kN�!p����)�.2�;WS^���@F�qQp�[��d�|Ч֌��� ���s��G�Nlg��ivvZX5%�E�s���y�r��B�d�E�n�o^��k�$�˽Μ~�gt���Na�i�[[_�ZtFŇo�O\��G��C��L���`���[�<�8
	r�>�)y�Ku��/P?ܒ[wˈ��#V�����Xk��k���K�nw�H>2�z�G�9U3}��{f�����z��!w����+ ��ZrT����#���{��a�U^��QF�t�K�?��2�	و��0W;�p�]g?Q�B�kNC�1aX&_�w�A5U�` �[��~��iô�{��j�
A*������/���[�tWm���4�<-��q��\�dE:����جHO��s�<����9�S��T�$v�E�4�5O^������na�;�%�Qi�F�ho ���3�U����$����ghI�%,ti�c��p�'�t*s4��G�A�I�}f��Tg.�!�!.�B���'Hѓ�FV���������HD���y#�d�|w�CP���Z�>W4V�����ـ� Њ����?7���&����:���n_�;i�]1��YiK}�6J���q�����j�@�/����;�RS(\<�)�̇DA����n%?�����o 0x������G��N���`f(�	�ԏ���F)_����#�rm�'ʝU�iW�������=f��OT*[��k������ ��9�b��FH���rR֓����T��$��(u��J��r�����$�Pe�8��jv�1�l�!���"�o�M�ڲ2���CK��\]BqbauW߅$���U�5�d1�SB� �ǎ�����Bœ?p�.�5Y�����_����\�⃻�O��G��}9�p]�{ x��#��D�� ����L�M�h����hX<+�ء`<\,�Z������o9\�t<���P7���C�e��d����M�90�"�V,�L����\�Z�j��Rk��a����W��=���M���	�b-��M�Qô��a�᧘�98���S8n)8��P]�͐��-Ɔ�`��>uon�>~���ٗ��aK�U��ߢ���h�,7��ޤ�9Y�aCJs�ܳ�Q�u��'k��y� �l�+�\�����խA6T���̲J::Ժ�ÌA"��O+Ӓ�@���\F�����}N��հ��xU|��F����X��hr���Xｑ��x��|NAb2��c�$ᒎ�b��f�q.eR�}z4F>��խ���?�G�W�m ?T���bwYC]�;�c��>�]a�\��r���=��6�Գ��#I��%J���k��>}w�D���,�� ����ә^� �OD9ڃ1�+r<���P�-vD��S�����3��.��ϭ����&Z����HVd�ez8��)��M�)�*xS�/�|�0Yn��M>��E���_��q�\1f)�4�A�VHZ�j>8P,����__ej�SKu��&3���SQ�r��x3����Qm(?�瞔?d���L����l1�� <��ǅ�u@Q6��dڰzJ1vᙎ]c�i\o͆���s�X�-��g@<�����C�w}�B���8�6@�7�������Ȑ]���8J�GD�mT�\��v\�o��׎��	n~
P[N*���B���0�U���s�5@��J�cR|�#�33X*N��:�:q���o�`��a���g9�x;J�YŮ�*�c{q�V�e@���NV;�2Q���ҭn��4ww���_g�U}��臮*����Ӌ->���hy������>�i�NSް��*�.��'Cmtx��t6Ai[��K�j� "����p�ŋ�z��w�����`P����'��@ni^w�WA<�g1A�c���<���;�x��� �D0X�㽜��P/�J�[7q����Gү����A�g��Æ4-�Vc,@c~�i��`r�����Azѽ�W�k о�=��oOvح��.���N�4?^t*��}rՐ��4T:����%�Z�y#Z�
!BUH1��(�f�TU�����M�A��F�J�}�#E������u�x�(� q�L��F!z]��J%�5����݋�.��"o[K���qu��$�<!�� 	��bv��a�W2�L(fHa!7��M~���_ε+����4��;�C~�J�|*p�: �&A�Nqf��}�dL
{����Yǂ	t��IQxR.@7�����w�7=���=�J���\Y�����k=�L�t���0z�{/M[�A�X�����R�>�U'��b@����U}��SQ����Jq�ת(eW#Q�<�P�P�o�bd�T��C��J`n!�"���	T�(�}�������nc9�p�:Ƚ������N"�2�����+@�U�H�K�	��� ��=wlҢP��l#q��O;��s���}��KW��k�0嶣O�9�!�,��h@�>9��<_<�����M�-��V����#�&�?2+�<���*I�&��Q �F�����LD��3_J�Ɍg�9ߎ��RM� �2�>�9@�{xC��'x�_�^���7yv ����VUkӸ4T��17JD��4e���:n��S�0|�͂� J-zl��"QL��"���\�0ϸ�P�1�)�u�?�͂>��V--a0���X�=��� �C��������½���Y0�e+rW�9��������Q�#��zs���hV����)@�zIS
Z����U������C�ƱR��U�V9/�������@.��vr�f�˴+wl�BD��W��6�5�g�h���G�f����\܌#h�qpff;��gG�_W=�C���]��ŕ\�(��y�˂���X�q'Jeb#�.�\.���-�cƘQU�x
���Olh���]"�-dT �p��@ ��v!�6���^�8G�4�GDg��:�N w_k^9��j$��{&��sxīTP��p,����R�?�WS�4C��}���Ꭷ�f�E2��V`�U9h=�Ӏy��W2�/��n�Ri�_!�~��q��m��xb\�-n8�M�k}%_���7�b?,�l����sr��]d�������{N
�Y�U*�6Rf�1cS3j�7����b��s$��
� >^�K���$t�f�c}��LٮWeR\