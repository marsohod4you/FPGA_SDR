��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc��3@���;��̵*T���që �|c\
��`P��o]L̛�鿕Z[<eLl˭�W?�;���Xo����^����Z�<�F�g\CT���/4�Ǎ�@�����(�Lx)�EF}��N�QÑ�*�����Zf�ϏJV�E������V�M>؆1"��0}��{�ƽ�`G�%[�,s���>�ӹ*����ںA��j�'j��''$���F�Sy�,�v��i^ٜ��/f���.�n���WG_�kQ
-,�.UI��ۉ;��Y��ULCͷ�,lY{
��B���<�����N�CĖ�Y���3r�����M�Y�����c����s�^|/&��~1=���T��7*r��d� ��X�P��x�Ǒ�w8hp���戕���"�j*�A(�5���y}Y'�2.&�*�/��ܴo���Х�si��� �[������K�7�{��俉k)E�J�7����$�ѧ��Xp��&P�{�̢-�=���"������@ �젟�\����&g'�'�L��$j��Mh���tq�)�<��!�������K�b8ps���ˆ%�w��5���	@���P* �;���F�f�p�֋��TרÉ�i>*��,�m�_ 7�
3>;~���؅8������1�R�����#�-��?Ӂ�y=�%*�ܻ�v��6�`�Z#X3q� �����s_���t���j��3D��L�n�o�L/�� 9
�'|[�!jd>m���o�σV������'2�ȧ�1aK��/���l��yٗ��~�!Oi���C(�z 4���|?n�ʡ��6A�g����kO*��Em�+�6� p���7|a^����sGK��p����B3���Қ8�~$lÁ	BN�*���ʸҷ8=�J���c<C�Ǚ�0� ~)�ǲ�Os5� ��amB!��X�,[m]F�:,U$fX����ٹ{��	�K�-�ɱv*��1l��V!1ck�5i%\���j�/X�����b������$	H��D?G�R���C���2���L<�fU⒢TN�<���?�[Ǒ�@�$պ**L��u���N���ȼ����t�9T#I&�硑k/j �7Ѽ 9�a�ޜ1��|6?A`{}�}5
�*�a�t6����]L#��%Ԓ}h��J���B�.���9���҂/|�{��8+�O�(��K�U�!��^��ӳU�Df]����%�3�q������ZZ,�ٚ�l�n��H�󞋹QBE#��lDQ�F(����WՑ�f��ݨ��TE�q"
�
����]�pr����U�bV6��gx���I�xh�slYODխ@_o�/4�����L��I��rp��M�s!��C\�1s�tkQ��aw�������2	����N�FD|#�i�kb]Oya�L:Bd#��u^�CX��UH��55qY�d^�#�҈�[ί��&���.P�뱯��^���V�YB~7�Q9�XI�K��}���b0td4�gZ�=l�&C�B���G�� F�5/�z9�/�r����orC��Ո����8��tG�ܴYP���EA^����y+8�T�ks����*�5�����A���95��������t^�B.$ȋ����rHЂ��;:Ro�B�R	KЏ3x�tR.��rz)©J��j�`90������p|,Z�xJ �pGZ���+^��|�!E�@����,*еM�v����U]�-.4�$�N��C���l�>�������s� �r�0���";��g���.��n{��SM��fq���� �A'u�t�F�^{Sm&�����.�Bi���U`-~��TdbNN�* �CuE�Do&��"�V1M+�b8�M)�I���&fq8�\$`}�!|ImᙂsR>x>�⼣�ّu�|t����p�>��q,�:$�ؘm��ּ����2�gq�
i�M�L�\��	�R��Z=�]�Q�H)3�b�n��R�UV@�"�UX��%:4�R�l�6!���L���Pa�r�Bߣ�/��{��/�*���d�Wy`*M�b5�%����KcJ�C@|��cv�	�
���<
��v $\}y�V̷��h��@�&b�R9�&�rи����ͥ)�Ka���N����j���,?!�8fV����K��d(���m�Q�4qۻ�1 ��㸚|�6Vk��2��ֆ��NyQͣ��TL�z���O�CmFp�u
�oj]X7�/��N�@���8,�c�kk��u��EI��V��#:Za`����DZA`�
�I�� �ڏ�ct��G �8��况��>Lץ̈X�i�S)f�`s�tF�}a�` }q��E��E;6�'�	+�p��R�TG�����q+����I���$�:�]��H�V�XK=�F�ɗ�'1��7�!�s�G���ܭ��L>'֦
A����\�]½{�jC	o��Vl=0�-[�2mo�YB�-M]`�[�J�=��4������t~� 7�$��Â6����[��n�q�_�(���L>���:�.aB�Q�C"P�ϻ��\R	�yu𣔓���=7�"gA���4��w�$�t��:k��9��*3��˞h	N�z翉u� �7yډJ��w��N���6��W���X��J�V���e=�-@s�Uq�}�\Q� ��+�U�qN�cȓ�`|"%u�	F�A���$��tu��6^�}��ʦ��M��Ϥ�T�&�'ق-�T���O��l2��.��[�`?t1؟@lv��t�05�r���gWt�����4��X؄�6r9B�l�'X
%�ۖ s>D�l9�0��;
Xx���Jv�˝2��Y�h#"�U2O�a�/��^��7i� �^Z��X�J�?�}�����?���&r�;ޛ?����i�m�zKX�.{\�b�p,2���;��ޭn�u�y�K�6�h��djh��im��C��5����J8r�w?΃Z��8&U��Yă0c�3T^E+���Uk��Tc`;,