��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��l_����b�-Vț�UM0�JK �73�h�J��ŝ��ܽzAV���.�z�POifK₿7�\���"q�������.p�<H'�=����B���=��t�����!�����\>a!�Vt��@#uG9��P�r�i�ʒ���u�^��/����c/���$�9>+�ņ�Z;t�O��aՠ;�����ȘH+o�E�Rw�ƮO)"e�2���3v<�D��O2?������f��ĸA@�EA��t\�E�-�"(Iq%0!BS��rYb!�~�����C�%e��H��Y=�����/��r�SA=�D' v��nZ�T�y/�-A���B��&��C����K0"�����ZR�k�ԁ�VΗK�i۞(�?�KQ�4 Vr�}� �&��n����M�`�=�"_��A�oaz�F|z$�A {����^��3���U�3VE�\u������qgS�Ԉo [�G#��r���k"����H�"�H�����6e|b�L���i�ψR��hmν0*o�2xR��ky+�6������><�):+�<(K=�+p3G���M���o��]�ঃ˃r�i�̱G#=�[M� 6��`xz4�1����ׁ���t�ta�t�;�~3���#>$�%�$�P�`�����T[�ˁ���2�;$�!я�y�_k�3dA8�2i�B=�M���G?�E��-V� q�rDjh�	�b:�m}]`��7�D8�
L�q��ir�ø�>i 1q'�N�l�_E�)��h8&4�U^:f8�D}	��Щ}<^�.^1"/���O��f�,��Ā��['�Āů��A�54p�v�(����TL�R9пD�
�DY�� 5cz����2���K��J2!X��ERaف�𪰎����Ctݎ��|�&%�!;�׀8'}C�P��6 o�x����8]�1�ŊHy� ����E�eB8��vXU�[f�dPE>�VY�)�y�LDj�􉛜��G;�Z�2�:����!���ȏ^���z�v\�~�~�0�1����e`��*ƀ:S���:����G_].B&����]���0�2��~��� �@������W�590�OX�d���/�4
�Ը�zu�m`��0�75 �� j��%1��9��铘���E9����q�/�0c����4(��T�۟Ϥ;x�*L���L��7hc�0֓��x�����{�)W0�x��jN��$����i-a�m�4f"�y2�'!�}mE��6�PKآt���Up.�(�6Y}��G���j=1�g���M���۠����-�I�{Jl���wxa�5� h, ;����eS��a��E$n��i�� ��J�e�{g��@=[`�.u�+���t��<�� sz�y"��><�wB<��CI>�B��s�W�sX*��H��څk;�]��+����m�E��(�rԍ���Ei�Z��Ƈ[&�L�0�.��O��	.����.�nk[1��!�	J^[��{�t�F�q���`��?Y��W��
�ʅ:��^�u@�9IvEG�K��f������$�w}��ė���{�Z�=��������Lr����[?�0�b�3�������.�J�'� ��2!U|�Rţ�cF�xT+��>�l;[�M;�����z1+�o��z��#����}ٜ���gw���Ք�VcT�U>R�}�`��y���4Ezp�d��l��OV�9ĩ`cA����Ym�I- '���BEKF�y�0�_�{:=�>*~U��e9�( ��p�J�������K뾜�O�\pg��c�d���U��k��u�!����Jź���� �=������#��j���Lc;��O���U볝�)}3j\'�Ѥ[me8�<ǎ"�8�	�l�/�ֻ��]d-�l�i@Uf�I�;R D�X�QH*�����keG����o��Ie�+��N��[���0��x���xB��> �_%�1������#U��O/��TTM�LkI�����Z��z�S�o5����=1��+��"8�ʠ�0uG+
y��)�j���� ]��'BҦy,p� �_X|�܄o�5��u�]������3�&�F�_C,)�Z8�VT6�;�&��_�Ӱ3������Q%J�
Q�o���Z|$N���+�b�Eqa��B-03jI�jRGO/�8��+Fm���Y=+ʎ�
�=���cE�̷Ld's.(�Y!�.t���Ym'IOĩ^A��n/y�\���w� �h�Ԅ6YLn7�r�,T���i�G�<�B�7�k��`Hn�������	4�e�g�����*hh���%S"_r���?t���Pkz�B��q���������Vj	��1���Tr�P��h�0�L��霁(3V�f�t_*ڏ]x\�J�:������������/o��M,���>*u��1^�n	k���0�#fU9NR�>�1q�ɐ�H�!\�� �n�8�H�C������֑$0�P4oBK����:�l��$�N�t����wu�4�;C��hɿ�Y�ӛ�2��f�#!�/��Ç�!���1��������ov����m�}�������&[�}_$�����nz�b��M!�h��H���@;����C9�H��z��>�,�.�|�l�C�cE�����Hf�'�12�����%�|F�H�nm�{[�Կ0������Rh��EӐ�x� `>�=X=r���g����ݵ���3*����h�[��Ūαo��Ǟ{��q�?�����n0`4�� �����E�]�a/�Vo߅�M=eMtw$�;��H5�uO�l����p�ߩ�I�-���X` d4r+>�_3܂z�{Z���%=4&2����L������F9��^$透}����C/��Ef�T"k��&!#3F�+N	RXAј�����}]&��d�V���9̖S7a9���[���xO��Sh�9r���j�l>䣊���X܉FL������ �f��._�w��F�[���d�9ՁQm�4q����`���>N��ǜ?uڡ!Z�K����#JFF�p��g@]q\�Ik�\�2N�������3���݁�vS��������~[��oľ0y�˟���_ĉ`dz[�!
�*ʌ��3gH;/e��'������U�$��S�Y�8m���G,ٯ�C()V�?q<"�:��O�0L� L������.m��ˍ����m�����s�.�0�f�*뺶��mȜ�$���z��!D���SF ��kPȗ.zFB5>��5eDj:�B;����%m��D�`��8�	��'\�U����}� �:���lr� �H~�8�,�")Z l�Z��?<�y#������'�"��mH7�y�3�D������4)=�`�ˁ<B�����gQO���$>�����
aZ9t:���&��4�0u���#o�82Pg�	�xj���И\��;�r��fA��8�c�:N��'d(Q�F�C����<�*V�V7�h�|����QO�Ɓ,5ù�tx���yeC�!H����n�y��{9lBf,K�٘þ-�� �F7�#𘌅� �}[�������6�ȹ�R�����\@��R}�.�J݇R�iLC�K�N�A�����6V{}r��%y.�����1.3�MTvZ�@�9��ͫ�}{�\1�aNHo���z�`2>]2*��H���[�{��ۅ�����R��M0�~��3���n>*�9]�)�
z	X	�4�{o�'�mg��½��Z<�HV_t(�Tp�paHF�%J��δ"�U\����Èʲ�y`x�M{�E�6�fJs�2 W��惁�����㊳����.����I+��h���Z�a����N���0�U����5 ���yY�\&��6�Պ��� �P(>��;!`�΅�.�M.����i���)�8xW^���~���,��x��#����ݰ�ŉG�J�n�f���g��9��Y��r~u"��6���w�NN� <�Z�1��n-�������#���GMߨ�`?�HT'�m�;~���y�d�G��%�=�52��,�Lv�8A�i/C���6<ĵ����o!�n��Y�g�KU*Oc�`0!��"&�ǖ��kv�"pF�� �Rm�cu��# �5�t�A�
��C,��e�:�+_�s�@�F����9��a�%�sh����Y�E�u�1yw�H�Hw��ߝh2�Pa����]u�?��}T��2"��B�zM\����}��<�3��e��(�8
��l�e<�59�~�/�?aJ���>H����5~GE���:� WS9�hI@�x���:����!���Ż*�?8�ظ��5� �!kJ�IhJV��/ xy� ���`ӭfԕc�+L[i8���8F�n�^2�悪ëN�n�
�~��f"��]������:�<��Ǟ��
��_G"ͽ�u:�v�=R