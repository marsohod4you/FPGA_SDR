��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\���X�Q鯠9ƚ�M�b9�M�Q�z�n�j���أf�W`��;ɿ�T�y�W�u��1}��������0�T�u6�&�m(��B�%!�2��{N�N�#&�3��r�83�v�W��V�_X�7	"���U|E�E�Fj#\�HD1]�|(�צܨ v|����nG.��g]���C�9[W��(g����8!$�[���"��5�l��ƨ��5T�����7�� ��X6~,ww�SY���{�B��Zf�pO�	����P'6��bC�gunꓰ`�Dˈ�p2���x�,9�"V� �,E�^g�ΐ�β}I%ķ8�ز2,��5�$� B]��gv�r/,�-�⵺@�G;c�SY\�����'i_���D�$|@����$ L���+�Q�XKD����~�������x�^dѵ���T�E���%-d��=)%��HRh�F���:���TNݠ��Vx>v9���>�-m�}3a�2�g�SaK��%q$`-�}�O|��J�5�2��D�È�ц`�����=b��=4�{��v�0K��_�����>#ƴ���t���'_�n`�K�A�0�O��H�`v�1Τ�J����▖p�I"P��������(XyEzS��9��.-Li�;��ۿf�nv��.�_�%}-�|a� ��H	{���˦�}%U��UwOWq_�R���P砀��Q��H�ºL�{�k��K�LLE>����ei3�I �)3�;����Ny�/���������o�e�d�I�^G�OD
ȣ�a)#mLUXk]_��Qj�]��1��2��V6� .<�v\�SU/ؐ��ڴ�7]gO0��������8�b1�JKk�"޿�H��ɯ'߃�O���(f=��"�N�Cذ���	[K�X$kķ�F�~�R+���� n�����pP� �L���yC��g�C쓜��#ɺ�����Og�H��0"��O��RK'�G�?��e�BV�me���Q��(a �[_����*4(�iM�h�38��zjۼ�]��^���C��2���.:������V;C��v�������>cydW�di�"�u��;�`�]�J��J�3=},Ga$�͵R�2�����WA	�\���o���D���D���p���l��r�ے���/�]�߄��,@.p��t����~z��A˾���C��˕`s��l�xp��ے� y�W��x��6�Q���m���oϲ˝]���C�=�9'���cJ��#��M 㶬��N�P�ߍ�0���a%a��S��5f4O��uA�R���t���t�?���0���VI��^?Jk�A��L�4��3[K��u�j8�fS@Sa�,���[R'�C W�])q7za�b��aʛ��5QYF���n̈H�	bV�m����-��K����n������[�4����"�IE��*��m�Hp�T@�`q�w�܌��a���)�6��A6qt\8[�L�֮�}��kx9
�E��%��#�9�OT�������V�W �1g��0]W�1D:%�%T}/���*G�0��6�V��5N�J@˯��z���g����=�F���ܯo�qz+H�+	��MÊ�R\+��9�i
��]��"�nAB�b�7`x�h�
w9�U���Q�|]��f��s �ۋX�W=�Wmd�kkA��`��IC��ѣ��-�|�Ď�i.l2�,(��R��;���|�vx�R~8��(!��A"w,���k6
������^��O6� �]^��%6���++pm�g�/;�d�J�4�v1��� �9TwA��f�b�C�� \]AP5�G\(�dy}��,ZR;�E>{C\'���; �\gg�(����Br:�
T}%����g��澔BD5��s��u�#j�ORV���y20,4h��uz��?�&�xN��N�9�^.����A�%��ݽ|�G;�Ƈmfu��nfQ��>���S��W���E#D�1s'L
��J3�*_�<��R�6�ښ9i}��7k�ii�{��$F�g^��PcA���Ȥ��Lg0ъ4�J�f�X ߻��k!X�W��_�u�\W�3fK-��҃9��������Cw�[���|��WA#�%��c�5+R�UH��y�ǐ�Z
Xl�#�懐g�?QZ�Niv��ײ1�I�a׎eP�ث��wf�$xpV����	�◿��ĂORμZ���6$YiN����k�ުD�~�>�`�����BC���0���$���x�R�#AtO���H�����®ٖ{�"欔�a�.����\�����6uE���������H�[�W��.|c��"P�U'!d`�@Y����a���ܘG��8m��	�� W�<�b�׆�W�sl�a�{��d`S�d�{�D:��O��Ν�7KH�ۄ]�y�:�4��N�Z� ZP
8�w��ʇ�a-�P����i�X��Y[�����6X�zzNV�uǁdc1!'��%��N�Ϊ㹹Bj��t������&���eͰ����Ơ����"���l���brms˶+��G0���:>��&���T��y�����'	����.PZv�d�J�\�&��\��qE%^�,�������W1�����X��&S�d�2�(����#$��l؈ �����^�S%��=�1���cƿ�<�1��r�x��+������/ͬ��f�����6�������̸bt�U��:�n��ӌIb�X��!I3'��r�ԳEN�X�	"��0`%�)2d hL��nd��G\BX�#����;;K$4"E��ʋ�\C?!����[���6��u�[��R��}s�A����-��B�'~�,d ���������o��cП�p�:�)�a�)Dh�l������V�(��6Mĕ��r��XzKru#λ�r�1Ч���u�-���阃#I7cP�g�f����l��F��k�P�%(&�_�w����Ldm_�s��! �Ox��qag�����K /��ո���r�LǷ��FUF�M�lF�]�noM�Ѿ`q�z+G�E���Uss	ÿ��"_�;�
�NiitԐ���o������yo�wY�_�N�YM\%#�>@��a�����)g%�,�1�7M7�KH�����.^���z�e��"+`@���A��14�a:�9�a��M�=]���e3_T�d���}"�s�h�y1`1≳�{m��u%�D�y|�aWٜ�F��7�
�>;����	���H;�'��8�ʈ�N"olِ�)��N�6�	8u��#���Rj����ŕ�~�)5���!��ȼXQ��u��s�|���y���@F�Z�C1� @F3����݂@���f;��D0ҏ�d&u���Ni�<j��R!�[=U��C�q�`�jDOt��@��V;�����9A�}n�E�A/��0lk�m%�+������[��o�,�=S�N.#s��:2t��fD1��L���V��=L��?^���ȩc%��B7D���Ұ*w�b�ԓ@q/P�)Xj�e�P��eJ�0Y��o�7�����WqP�cG&���]P��.�`wS� s����xK�'#�j���bK��tbB���u�.�����u�� 4���s��`�l�d�4q�G��g�*N!�1�p�FVV���mK�����p+��튻 ���B�d�71r{D+�0�����|4�cCW��$a��ί|�����X�Q��܀ew1� ����8�п���A[PB�NCAD[��F�I�G:{6wT2u"�`�!a+��5�(D�,3$$�u�8K=��(�E*횏�OGl
���,R���Pڧ��_�Z+.�"��٫��M�Mf���t}^Zd�MHDt͞�~��,��������&�	�}�6�]���T��<��S���
.��+�Z��w�����qAIJ��ɿ`��sR1�D�O�lHAG<�G}�$զw�t���l�3(��7,Ne�C���mR�_�mc�&&-{:�ǎ��̧��7�"��BU�4pF:"$�ЏL�"��l��)��3���,(�=�s����9>!�3d���?�+�)N�|8��d��dU4N��
���M�`}��=�V׋:@�F�e��f�	���^��>W%A�,O2��G�Fx'�_7�ٕe����=�����>���Ƙ!.8H��3'7��\i��1I2�&/�1YWu� ��O�w�j}tt�ᩮ�]6p�R����q�)���D��o���ol�~�I�:��#$Ȉ�Qד�֑d�A�H��),��B8��i��`�v��q�ѩ�m� �D�N���f����\�Ϗ��&<�@���[T�]�=�~H�&Q�T����L^D	c�WM�Ň�n��O��GK�#m}�BA�oR��R.��m��k���!
�x�u�T0�4��:���jk�N��&�kn�[�xMm��,�d��1y���<'��&�������+�in��'������6��'��]Hv�/"s1_���s�[��C��K:vk�0�%M��딊ƌ�ڵ���̉a�?5z��*�Y�A�_�嘓�6�<�c;��[�ao�
w�we�*}XmY���|L�c�FL@qǊڤ` ���u׾�.�n��6�r*7�U[�`�˒(�W���Wx��.7g?��*�\��hw�D��`A��,y�p�cu�V�[�،/�+���������q��6�.{�b)��8��09�� ��0YqטY��bmbYĨ��J���#Y��MU�oW�����Y��	i�XJ�wg��"�U�G���"��N�"TQ����oU��V��뫄@3��0�[�f��"0�@y�<�U8�������F�@���8Y��O<�^�e�� �͈MjC�32R��	
�"mUK5���cI!n�kʙ�-J��
��#��P�H��S07�}=T�H9n���E~
���g-�B>�EK��R�Y����U�=�೒�O�GkW(_
�M�+�N�8 hF����W�ʤ6�k�;Zm�[�7%c�
��%����MZ��u���<×��aV���v�d�bmh��7�{:`��j;�&C���BGE� �W�U%�-i�8��F���Ƅ6	����bV�K������0|��__��k�@�ع E�&O���CuC��5��(c\�\!h�*�W"�` &,�����o+�������4(�:u���苣t'V�rݹ���0?�VV�l�-�\��s���Sk�N{g��ú���Ǌ���~�?}1�ٟ(�GA�nR}��f���?^�� �J?��L��/�m�!���F[�o;�p��vE:E[U�����2�oLX�a������*el�?i�K��T2�`��|*�_��`�k+�Α���9�G��k:�ȣ�0�D��U_�Q_� ����6(�Ytt��0����~�R�E�wٰv��@���<e�'1ʏ��RMj�'B�6�Z@�n���nm�%��I��4p��ޢz��THK� LZd& SL�)�^��~-ˎ�a��.�����6�c�p����O���G�T��Ϟ���(p.mP���H��l�,��������~VΧX8&��{�NP�HEqOB���k=����̢Ṋ �Ɣ>��I"��O��<Ow!\P9�Y�?%SC��(���MS�ǆ�`cDK�K�I@�7��A#58>��(�m�����.��>j��Q�yui7�6&=�.¨�(H85�&e�6^��mU����7�\��z�6&܂�49:o+a(��֣$�au:)�pL�Ҕe��/�� �f�-^���b�h#��Ƃ����F/���?�<��r(�ԗ�l��
l���Td�&�^ħ�|"T۠�D�k���NM�:+�G�ƚ��;Ӎ9W7y� �"�z&�1x��3�A��~V�j�l́ߤ�m����ָ]���O�@����!,~��)��!���smt�X�H'�OU��}Z?�ld����6Tm��NJa�mZ�H���H��¨�Y��/w ��S
Mn䄀�J�s%_[��5]���mt�RV�2 ��A�	���D�=�Z���/��12�}��\��n{r��̬���/#�-u~�\����zP;B�]�X��X��Ѵ0A��;�f���j�L0��<�5�B�s��]���{<k3��IDi��+:H�C�!�V�!�C��kwp�m&�Z���Epx5��q�M(`j�2�5f�mu��!^8jo��֦F���n\d���AH�� ��-=���D��bܘ��e�qϿ�y�B���m�q&	�._�(��2'�.��n�y���(�O��L��.�{�L������Z2BgC����IU�����F�ldW��`��X��y��[�m�s-�!9��1��픑}���!�!�X;oWQ��=<m;�mF��� ��IC�V�.��{��0�,�>�̪މ��b㓋s$�g��3l5U9�	4k��(������VE�P
0<:gc�A1J����9�xF��'�#�E��>w�!�ʬ��f�[�C�h�g��*���p$)E��T֧>�b5� ZPQY�Ы�\�Xr\(��]���+�U�
sX~/a<�'�$����"�S��U~�K��O[��-==,�,�P.@1ӊ�{PD@�6�&��2t��M¤j��+�y��{�b��Ψ�P�;��f�whA�	�$��yth5�d����9�9�^�s�sJ�� �(�� (gߺ5��I�8�@�l7��x�HK�Y<��r�du���=;��ɦE�]��@vٔ��9A]�**6��-�ȹ�����^�Z�(W�ES�c\j0�����I�s�"���K�9_IL�O>W���yRY���w�r��}�,oQ�ZE����nG�s+� �%q$������U	�%��{s1�W��KӖ&?1Ո��<P�a�Bx�T��z�̨y��F"xM>�e��p �E�+��"���Z���dFT|D�Td����\KA7��0Z����U�Š�f��nt{p��s�#�%3,2���kJGX/u�0qV3jgi>��c��=Q�Nl��J�N��HhA�y4�Ѓ�[s|a��ӈ3c$K�����)��+Pѡ�+j^�24�[ԡ�K\</� r�0w��)��k�P�W��oϔ���T�>��'[��q�-X�λ�=A��!Y;rӈ���ؖ�"�6{Y����r�K�QN�����}�f�7YJ�e�^���ΐ���|5K���ؼ�[!"(Y%�|@�Չ ޻.Xz5�$�XQNp���&�m�]���N�lf�����M��õ}־v|�A�`��C7Q�u0T���_�4�@UPRc���~�$������ĵ%>m�
X��.ۗ:��3I̾Œ�A
�I��	O�N�^p�L�np�_9�ݕKV�%�C.һ�95-t0��%�2.�h
�^�I�DUO�8W��յc�j���R.�<(G�_ݚ@Nw��84?BRaWp� 6jk�(W�.�6���C��A�%��鍊�ye)��$M.�ne�3��C]�X��3
O?S��M�~�LxR������hTή%P���#�vG���H�����$��I�k��SRTM{"���P�wGo+�kM:;YsE,��ȕ�m�ڑ�qù�r�����S�8��U��	7��������CT�s����*>]{��]��O'����F�4ިg�1�j�|N2�����"��:l���f[�R�\��/��<�|-�Z��gnex�"Ez|lzޔ;�)���KV���K�mfB���'��A�L�}�>r�^�����Vԍɀ�\���ֱ�����|���"^��{���P���ow'�
���)����2�$x�����[��FS$�k�e��m����.�fVC�[��ֲ;�r+��j�]OMn,�"��U��1�X�
q��ہ��ex˷ʔ;ň�%���U�_[�g��z�0�L���2��ݾ��_�I�l�_F�J��t怯�쳪]�v��f��WQ��������lp[.t�3�)��{aU�5z|�hm2s"�>��$��ɭ�� wX&9�����ô�*�	H���:��|��eI����r#���ߣ\��IR���C  �n������a��W�c�|aƼ!v��fŝ�4H5�7������=�U0��BvK.��:y�-��7�|�7 x�A�T%�D9+�D	s��B]����G��B�pQ��^
��.zn���%ˬ��`�MF��P&��M�/���0�����dY¦&*~�����	L����_����V�ܾO{��Z��H�>7�*D�[�Ȭ�}�\��+@f\U de�1=�x��: �G�%����Q�M�ҨVY8���5:f�����Vu��Z�Z^&�_0dl�����kS}<����;	�fsӸF�a�a���L�,//2G���F	 �}�x��me��N�C}��hp�A
��p���V���W<0)xn��L�v�/#{9��夗�05{�1��n�Y�wG�;��+qJ��� oz�l�ܱ~��Xɕ3	!�������K����%�@�~�x�L�0�Y�Zo�#v�\3s0ĎBG��GS�H5���Z߈'�J
ZjƦ)����	��X�B\L�1�UA�t!S��J���儚mS�NB0��) �0xۇ->:a����;�q�U�i����,����W�vl�Ԓ,ԣ/q�2ve�}�)�B(���n7+JZ��_cG�ĤT�,�I���Ma4�$5<YfMg�̪��^��F��:�/#��~a$���� k3������u.0Q�94����`t�Qr�x�zE[f�7[�J<�_���@0�U�Ff2�7g���N�U���5��p{��1A���S� ���\	�Q��:��,��>A�x�}��.δ52)쀙�j�&\�إ]kA\�d��n)�P���?���a.��ǰ����4"h/`�{�-sq9Z��W���포��5jaJ����+뇛�$��-`��b��#��v]�Y��x��5�bD���d��M,����{�n�1݌;$6������L�d��p����B���t0�k[7AkWrAܥ��7��З|�|8b�է[�.�1�ׇ}3�_K��3r������p���������I�	!��
�"�𦥖Ǆ�U�i��Q��P�N�Z$o:�D�@��i���'h#O�ժ�Cr���i�i>���T���+l����w���9�;`����]%�^��@���R����i���W>�>,k���6q��`��~#'�hä'lb�?� ���z��|6_GׂU��|>#�FKj8�#�W�P��T�t��\R�D(�g`[L�m hה<�兰H(�(��@�ٷ��|.ۇD�
�s�=�����
fk���sZ��C���Z�:��b�8	��]�]J�i��2S�*�s:�=�ev�g�d���wf��&=֮���p)hMe2yub�����s!S �Y���G����j�OB�,�yx7㿦]E �(�Վ���${��nd`$VzŰ�����#ੁ:�ֻiPC�ԣċ�l�����Bw�{��{��jU>�s���]���".w�$*I��,�>�ډ߱	��	K�]�v� ��{����s5갂�)_�.�ЗI������&�jI�Mo;r�\Z���ǖ^2�jv��:F�#��Wp_`]�ڸ���6p�S�+�����,cLǻF�P�a�xe�*��>[菪�y�>��yR~��a���~0��R_�r��B� P�Lwg��v����qQ�B^$*�-�R�ֺ�d���,3�ydQ0�74*�-i�L7,�,�)�g�i��Nq�xl�pI�H��l>��*�}���12���'�7�u
�{[��hys�<{6?v�G�h ����ٞ��ݜIZ<�:��f�tK�3��ۄ�Ys�,U�T���7P�@�0��횼bn6A���U�rz��Pk��F����>V#A1�.J������30��|�4��8����a��p�T�b��b�H���vs����d�dW?u����=xzjRe)vO�#�me۞]e���u���C��v�'Z�c��o`1��[g���m=.ݎH�);�H�6~[��s��֬����O�
$�HCⅮ�Fk{�RO'�7����=P`���J��/�h��*N��k�l9U����B���$/�r�,�n���7~�h�b�\m��0'�3~�έv;�q5�}�ir�^��G�dzV0.�0Cݢ8��K�6Z�`�h������I��R5��e|-&�����������0�+ê\ ���h-v����5s���kJ~=@��3�*ѽR`��l���2���J/J�Ԛ��!c"�کJ��Zi���i�&0(D���w.Ԛr�@����>�Sq�iS�In)LC��"?"1��-���쭯�I�z�!|97'0��[(�?	��ڇ'd��U�Є"��FP�<3�!Q+�:<D8�y�����4�*~�+�����7h�
�?P����8���=e�M������4'2]3G"����͞�h�d�[Efa�%���9�T� ���聍Xc���kc��1%룦zu�����1���8�:Sc�Gc�0�,�K��J��G{J5�dA�N���Z���������:P��u���ks��/�8��}������	.c)֢��&Q����	�����j��t"�۝��+���ޑش�gӋ������)�����1��ۑ9���	Z$M#u.���� �Y��F��!���Uf������YM-nȮƙ9�z�)�p�T�8�Z��ku�?^w�F�xvk@�29%�>��V5�:#	�1�R���֚S�T���Jֺ��۴�.�����1�ԙ�0��e�Yl����Nϛ�/~�
c�qlO(����ߢ�ۻ�q^?B=/{�e�4�)t�S�
D༧�W�x�3��x�;B��^�a.������ڼ�StxЄ�`>U���ȫ��E3qKڐl �쯻�,Xs��'��8�$��B��(Mt�����^}	�)��غ��17g�r�S/ja
�WK�/!X�s7���@�P:ۗ�[Ij�M��>�� �������WI�̝��ف�"��27���z��߿��UQ2G7[�/zGbO�]3sh���Jh��K�-�B�t@C+I}�|����m���|���%b5���:��<фhG{�b��"zr��n2��v���vv#�/�)�5)�k�A��q&�����_ߦ���X�����b��y����|l�b7~���N)XC��wQ�	�p�;�#Mz�Mp:p�>!py���ۻ�ܲ|�	z�M�f8'�~ ��ߨ���.�>p��֕~��	����"�B�d��d@�b2�f��_2���8g|\*$�a��y"G��5S"����bpU���&�l��-�6܊���6΍m�
����+5j���T�k~���eޛ�RΆ�EB��f���Nύ$�=����]�^ѕ�F���rn����J۰uAA\X�O�c�����o�%TLQ�V��B�4��lg��B��j榶$2���"��=����4�䥆M
7 I[o�zll ��"��?�.�;8�S��d1�A�cE�lM��DȥR3ت�d���)�F9Č�X�Ԧ�C#�4�Q�U	ā�C��m��������2i�B���?a+�}O�z�41��/�2�d$_Ω��R���k�z�W����}%�Q�1�����IR0�-���9*_��YT�˱	����u(���T�y#���v�h%��ᛦCL�����}���)����BmU>��+:��3JC�d��le2��=jғ�Q�[� �[N�B�W�r��a��i���^J0����l"�BO�����B]ؕ�lT��2#�� Z:���C�eD;�^ZZa���U<'�F-���+�ډ��?P���K��F:�0��uI�d�+E>Bf�o�����ۢ5|��iy����$�x?���l�3/zl���v��ݧ�ؘ~W��K�ER7���V���s l's �"�>n�I\���H��"muО���BQ"-�yA���4�h/���
��\��A	�kc����+�F��&p�HD�Y����W}���)���Ջ[t�MQ�֥t��Ѡ��L��^������h��-�̚X�+c��4��<{�$�ˡ�W"l�����@kT���{�Ÿ S�X����23� ��M7L�Q�Ii~���8X�K�_OUi�E<�����!�;�.���G2p�ɶ:[
�ܶxb�C�4�y�����7W�ZM8�L�����Ł�d�Y	>��ϵn�����ȓ��"�W3Gi%f��r\��d�K�-<�$y'��Y�ޅ��B�xFC�Y�.ROԯ���OMׯ�R��}�ݙ�2��l~�ܶc���ĭ�F�~�yE������e�Q�Z�5�x]���W���x��&��g�$d��mHf=s@�`r�av��<�)j?	���hrUDCdMP������G#j�d%�۬KZ��Y#V�:���x��1tJHG���CV\rôƧi˄�%��Ss2�R��=�.5]��d�3
2v�` k���i5�MyA�" �今��I�?�9��v�m!�۬|����y����-���r�M���Έw%�D��̳�Z���y�I8�7!�T'�í�^����c}fS��!���D2���^3�۩�
�d��l�B
D���tID��iS�(��D�|z�B�ŷi�;2���ݾ%�	�`D�kMx@�_Pu�v�W'��A3(�ʑ"ۘ�/mb�V�0Ŵq���`�� #�:��Pt�)Eװs���̌�]���F�	�	�v9�l�4Ca�G8�`u�B�C�{� �R��-֙_y˫udfr���F��o� z�#�����k]��H�� %��Go\aa5�d[ѐ�$&���ՊUz�2C�4�� ��{@A ��E	�Q|u ��� x)L��F��(D����tI^�u#�X3G�C��O��F���(�Ftk��P���޲���7��)a%�h��h�X*���T]�
p
?�^��m6��w�%g$��՘!��|�h�L��8	I��fD�y�V�m����+���]FQ^/8N��E������]�M� �S9�}u��Q�Sˮ��o։.M!��ɩ�9"p�+k.��0ޖe�ɕ��or�\�P��N�����'}L2.^;��c�F��/��Ǥ���9�D�3U{ω��6�85M�[U�d�V�o�*Yc�3�NN=B�����M����"6Ll�3Ar�����<ο��Xg���M��g7SI9�h���.��%����n3�a�,�t+�Q%�����!��-�7D���܉�/�N��M���l�i�̬]�8hY��&KF���z�>�>kP�q�J��F��y�Ҙ��s�t�QO���F"7�	����En������0g`�/�aT[�f�s���7�1�P����ziߓiy��-=�'"z����ЯJX���S~8�U�yg�v��K5 �AY�>T�$���<\��6�qc�Z�Ɍ͈,�4�T+<��=�c��A�^oC:���O�1�[�ƠM2c
���:�&�uG�^A���Gb��3q�gm��B�E)`�c	��@�
x���uG��V���g�L�ޮY4?pњf5�I��J�!�*�rʾJ8[}�[�LL:�|e4Ӵ`0&Zc8@�ő��@�}RXHM�����J�W@�`���b6&:!/���� �H�R����U&�l�t�"+�i��l��xV���FmC�Ҧ�Z�i�UB�A��`+�Z����k�WZ��0���:c�"��/��g�b���r�S��7~��c)���lE�~!��a����HTȞ;o,�Ő#���XO^��Ew�\n{�B�I�p+����>P�/Ll��Y^̑g�pm� >�4e�a �$!�l�F�{e�'�N�!+Y*�
�)�L��G�6��X����lgA8I��q}`s8�d���-vdd�0⡇�r�w�V��ZM_���+}=@��ah�Y����)�9Ovk]��u?I�@'�&{�3��GRMP�4�������_�u��zL�0'��2o�8sG%0V�brǻ
�Xn�mRc��S	I|p�?��%J2O	K;wt[w�!�}F����k�����N|�s*TeKLD�?���8(>�����N%M�MӚј5LY�h���`��l�_(�E'��J��[%Qֶ3��_��0�Rj��%bN-����8�?����ל��&�Mњ+�x�`˞�L�1��ZL��{�f`� ��s�J��S3��4��՝e�����y����~|g9^�$���7��y:��X�������X�9D�i�-�<��:��.�1̠��-�pN��T�����F��/Bk�D� �8��]�P��e�$��ovA��5w2�u7��W~c���+g˳g�s�����HI���3�"Ӝ���#!c��+7#Rr�r���-IOCC(Z���Q��-Ƨ��Op
����'p�K��ۀ��0�F+��{��? ��]J�E��Q�R=��c�u�ĉ_�|`�j��@�U(��o; ǢO�N���	��$O�x]��&k+�Ʀ:��!}13�s�[UB,OA�5�y����rÞg���\e�8H����Y�3������]y��aVL(�����	�!�e��ɱ9���O����6�����7����y�N����K�tcu��zhr�A4�_q�'Ǿy��Y�3]�bˑ+�����v�<%A"�� h��\����|(B;-Q�������߂�^�<�5=�^�W���vi�����M��d�cD5:���#�fT����f2�P��a��,��r�O�������j�?,�n��&�+�h�����_c���k�G���q�{k����ycP����0������i�PS`^�p�q��ӌ?��P။/8I患!�x��#�(Wq���3�ہT���l�xI�56��x,%�}��_���=��ro�[I��o�B�*#%W/��^f���y��(XP�'�w�k��.�z��q���xH�V^Ӱ�i����\6����ţ��s�$(��@<�yE���oY�TD���r����~Ƕ�I�5ÊZ2,��<KE�%����q�=	�7���6��r�:�,@�i�\ݪ6����ѩ`OA�2}�V��G�%����W~�������%��]�C�=d�"V����9�/m��:�T��� ��n��s�5���	|�~�"�&A}�[N�'l�z�%���3=VBz{&x�Q:��KE9��»yj�r�c/zح0z6b0�n⒪[�����)ԭ��}l��;��Bﲞ���Vl�2c-�����}%oQ���c�-��v'gX6w���'w<�ʨag6"���+�po����o�t������È?�4��k��I�^&�uNj�ސ��Ɓ�3c6Lxk�/�n]J��`��X:��OR���]p����F:�U��-�%U\�|u,�E�g��>ԣ|����S�=��{�(��x��$ݔ�O<MR�=���:�u�������7�Қ��ŏ�Y%)I��5�_5����O����iyQ!#�*� M,���W��G��I�[UTI\�c�}XMe�=�GPl;��1@]u0���x����2L�BZ ��ޤ�>,��OIB��r\��ҷgG;D�<�`I��o*Aے�~���h�ӧ|멽63�L ��Bt�m�:r6� �BZ 'A�S0[�D�p��1A�a(�"U��/��,%�Oj�F�ܿ�jFc^�-cݗf����YʫU6s �4��2[�yP����� ��m+ʗbE_�mT�����f�B��3iqkj�k!�A��"s�53NW���#>��E���x憴�ٗ�Q��Ѝ�ǆ��L2ݘ�Pha���n�G)J��7�t�:'Տ���օ���T�(��<ݵ�o�����R�l|]����3z&T��[�3��ع���9�&O�dKK�tc��^�n��s�X-� ���E�ς�؊��F7I$��rYS���N�l��x�ٝ�Lv��d��C^��w,�\�R2m�2E�/Uq�@De�O-.�� ��V;�����/�2���������eF�@�B� �r�.������T�����"\Fu��:N��*Zcry<^��s�
!��
��<�Z�֢R
7g���4u;������/6�Z#.��/�EvMf��vc�ĕi�<�
b�ͫ�P&YS�4�T�o���Y�97(�~)��#~~��e ٩Ym���I}z���X��>B�]ӠZ)�� l��[��&~78�2��lΐsǑnڬ�z��M���4��os��'�:4%ʍ������z��7t��6�נ���d��~����P?��/���Y4�m�XY8����[d�jMQ���4!��G1eՀ�9k_���jP.���u�v�Pk#��s��<��������?y���-�qM����!܋\��'Pg��o�5��D1�z����A.�W���5��wl^Ծ������K�6��N�:�MXg����q����/�S��}m��n�.�@��{�bӜ��n���c�kIf��/3nu2���u�] ������b�x�m�C�'m'�����;�V{/ȱ���A52�z3�!k��F�X/��~$�kF�P�N��^s��0G�	�m~i�����S��}ߘ�M�܇��R���f�s=N�+e��k,�V�ν� ��3�7�b6ܞu݊�v6�U-j��f>�j,:-u;X���|U�5��=��nH�Y$z]��N��W6dȺp[��`���p)pmc  !!�'U�����#��s��U�ݲx���U����%��l��z����(;#������Y���14 ��ЛH!8�O�w�qLg�G��ė�1���lXDװ�9�#�P��:A#K �*�B�k��OUjK�S�=u���|�����@+����N�St��h��S�'������1�eѪN��������$��\ՑZa`4�������ٹ���ֿ�%��jjoPn�t��Ͻj�D���u~��sv��#�d�E�=��Sy��?��:�N�e_�{���(�k��xEF�����d�tmo� &�6��p�ew�5;���^9(�Oȇه������-u�0akhHZE�$�tZ����$��ݽ;M�]'t�q�U��mSq���eK,����8\`Mznu�fU�l`�@�ɭ|�sgV��G���(}j��g�,��)YoG�쌡�'��so�5V�"���������6;Za���1L���F���ʪ�^�~�B�Q��x�� u\4�>�B��Vz�8/Ѥ�j�˚�"vF�gj���1پf9���&�K���ӲIn����A����?K��3}��B3��x�S�a����0�\��������w�8������('vxl-o�w���NVm�jp����"��W�V`�&��_��+r�D��sq�?t��6f.v��F�Z�F0CHl�7�ٟK��.�o����<��a�%�<`ؗ��d�au�i�H*^)���tP��>?>)��nO+��^9������\��X�"^�j�R9�0D���$Dq��0�Kd�%� 5n�����EJAiu�![��Sfa������Z�O���m;�у�v`i�MC��Aޮ�	��`!N�s���ą��%wD�/��|Y�-J��W��|��"g+�HR�+�$�|B|�p�=޶�����'������E�L�|;�\�����Lnt�g��?y�8]�8���ft�� ~��&��-�m����;�����7�����G����R��&��_����Jf���1Ҙω�˙4��e'_!*)9�����72c
��E(G�ֿ�ӗ�����4�ʽH?���^Ul��(��������wy:?��|�ON���_������?�Í��7�C�V@�F'/c{�F�l.(��9���x�gCӒ��������F��ō�c�o��x�e�u�|O`6��c��kƥ'��_��<�f��l���f��xi�����30�5&�H���GbF0��������m����6i�y�\պ��� �Y[��oG�K�����Z>қ����^���t���Br�D�$4�p���&1��E�<�Lx�~��|o�I>�zU�|�~ΩN�Jb�̒��]�Yu�1Y
��wca�K(} G�j	=�gnF����s'��G�mFb��^��y�8~��Zu��v��2q@g���i����<-ĨAl�=Q�gBʦ��ȗz��\�����m�L�x��ޅ�"4M��:i�����Z(`N5M�߻�efc12�yoQ��O�jqN7B�<����F�}y�b%��f�f��Ԧ��@ϾB켒��5� ��P;�s���/�}�������z]�����_��o�#)lޱ����>�dȫ���aG^D����cJ`���UTgά#��S�<ɂ|:����w(���l�g�>���^�N�S�N��g��P�4V�[5í,ݸi
^��C������ϳxӞZmt���舭l����~�����U��P����N��#��(FF�|��a��0K�e����bs�r��@�.E����P£(�����P�A��C%�z�~��
p�}�{��}������|�M�RH��t��ȖD� ����2�f`��_�:W�K�o�\Y���k�	`ɬ	=���������d�:�g5cT�!?R�K%�?Mb����ș��a0:Z�fW��m�A���kƃ�
TwA��SB6���L��8ד9��MN��VZ��6Ɉ��)�W!/$t�V�a�^��}i�Y�G��η�g2�oM0,�tj�kw�g6}�O�r!��f�48+���k簾p�D^�EB˳ܲmr �lM3�L.�mb�$l����	I�����]R���3����a�Q�L���d�M�W�g)Y~�5�1��<@�f�8��2�0���}͝a9�M����R�¤�] 1�S��y,i�,I�\hb�"�_����m�(�h�2��n(k���(g��JWU��)m 88��(���SU��{�8���?�6-�����yog&@�7^���bE�;�=����#�D��A����w�:~6>|d&`���3'jM��
��f`�0�������D���B&_��=ep�~C��A��v����K���/�8�X�Ҷ�+�\�D�_(x`��K��,6;�U�]����G0Ȣ<^_�������r���զ�ٙ�B;������?Ȯ|�33�P���W:��*7������@��B��m>)'�VP���$1u4W�o.F-�x{�rg��`RiY'�,-�U��U{En����0F���7���S�>�Ţo\�����󆫌���Š�$L��(������'��F"t��g�&�%�pt���Q�|9�M���@x"����P��`���x'������=�]�'���3��N��ܲ��]d�k��ω_?�) ��WOb��=���
Jx��x�ƤEK!�0:�[����7������l՞+^�w�>�%B��=�Cn�0P��T��o�{��#��r��(�Q���r��7�o~�f�	ktGŠb�����u��!:َ��*���Y!���]�0�4�v�ah�󝨞�WRu?����\�Dp�)�w��,.��f(��xEH�l:yf鼗��+I�<Gѯ��B<*���6�F�̾��y���n�oYI82��� >���=fe�sYdGS�q^��a�C22�lc/���h����K�������7&�=��{�=, <��@�%0�8=���E�'��ʉr�h���R{^+9UF�h�|�q��'�Bn�*#�\�ӆ��3��� �������)��R�2+}�<�r������u�e��I)��L!��F��෌�^��D@4I��� �v�����aWz}��#\G 9���n�ү8s��7bє�E�ȃE��-̌���!B�q������+��QDg_#�z'i���ը!
�|�[9���m�9۽�`%�����e�����)���X
DYGL[PG`6�,�(��4�����E�!����!j�XH���9_6b���v�*�����<R�(ݟdy�a���OA�ؚJc&"�R��An��v�H��Q8�N!�	~�ʪ��}hF�gJI�R�/u߰.8��:�D����6K4���J�2�R�`��*o��,&��'��nm��:y�s>;j� ]��F�m�r^
��mqէ(�~�8��a�1�}��P�P��z֝oj�����2�;��Ib�?-�{�t�W�Nt��H�b�\�+�I]/4��9p��zFO�y��~��9�իg_�p���qT�=���=��e�������vM|9� �Y�w�!	��d�f�Fq���Ͷl��}Ѫ��F����FmAF�fݧ^�g�_˂�4h����4� O�r*�A��vd��z{� W,24эć��Y9��0�D��{�My��j<.�gIb��t��KK�����^d�QS/�����u�9�KhYR�I��.�tҥ��y��j
P�CrjI��	)z�*��z�HnF|����c�k6ueB��g�9C=Q���P�!l=f����0�R+�7��a=�P�M�Jb_B_���B���"��O�F �����s63,�Os�c�QB}�`�Yʙ�\J��W@�aK�ژ����5JXDߜ�ߞQ&vhPfݏ����|&��yn�T`<�7¿Hĭ���Ws�6�1��'�c~�I�-��$��`����
�jf�I˘$��p �d-�$�g���A�;���X"� �a?3�e7�
<$qUڪ�[)��N��L���/�;&��f�j��6�7œ	;����M<x�gas�L
�@���
C��+DH
`M�Y�?��� �.9�ys�����@�gW�������왋-�Z��1���gd�O��RX�q��w܉eA,�YR�C}vl z�+���S��\A�c��{A�ijy�Cr�Q�$EE۪�j%�λr�9X�������3�Ҧ����d���M
��)_cf��X��b��'o$���.碦4����N�X2ӿf0�=��S0� 2<��\���&5s0˂�C��ϛ��4� 'U�V?U
ؓ���̄��L$ux��Y
O�o�?���/aH+�fDj�"i������{�R�ic�<͎6�|~�u@�]m0�����)�V���yc��l���NV�k�*7�0%�+U;�m��-V4�_��^w�I�=k�Kur9q��[�62e˪��i�Ho Ub�zG��C8��������K"�=�;�C�A��� /�ڈ�b%B�L�����3��UNhJ���s���u�&��ց�f�Ǳqy 2k�,��Iím��J|��T��򬴘��i�
<@N�����׫���F��-��	����*}9��n��J="�I���A/]��M2����9U6�H����2��7,����,7Ŝ���^�"�k�z�n�{��JnF��y6��R��1���w"�k����ua�6�u��C��ā�}3��tB��o5�� �L	J�a��ѥS6�OPצv�Y��~)-�A����l��ئ5�W���c&�J0���ԽKC�g��bA�M�ҷ�#�&�����/&�o)���a��j�`JPK�x�(]���O6�6Z��Y4O���� jQJm�f/3H��P�2�{P,��uK���O��?.��喍�Y�r�=ܿ��.yoB_�:�F ���(ѳ�rG�E�Sb���J)>�rU����?Ԓ�]���0}�S�詀>�1$W��c&�rU]�KCo�� -���B.��{�Gw9��
������,Da����h���8 g<x�g�a�|/'v�6�g��uR�a�K�އH���"C���;Ȏ`]�����	��oi����s7�#���OBC°�S�w͞`4�O��aݤ��'Є�C��ӢF�~����^�tHz_ʣ�_�Z'Q��W�y���I�P���c��	�Mo�î���'/���0j�A���s����]�Ϥ8���y�q�m#�0Kn�����e 7�%�cF����Ϫ�����.�o0TB��)c����6SQ0,S�Sc��*�r<��Ȧn��X�.\*��5{|ٗ1Ԅ��@� ��yy�~E�j@УqY,Զ��L�l����/K���|� ��>�\����R���0:�ʾ��&=�!��u5O�{[_^�	