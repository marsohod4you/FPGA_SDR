��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>Q�y�`�}Cj�L��#]x�9�Ժ�-8w������G1n��� ��z9(�
jr�(-� 5O�`��K��P�=�GZ�L��#B����)��l��j$p�j{u9��7���R�qE�VfY�P�(�/ؚ�{
��.9��Mۜ�/ *�\ā�x3�?�׃��F�����;��4&D��+�{��K ����,hy�#d�~��,ePr�=˝a�v�o�lS�@љ���qzz7y������"D���!՟�aI�F���v?5�����D(5�5�Cv��'E� ^��b���XEtd̎�j���0pό�Xh1�@��>7$x�U��"(2ly����#t�i�״$��K�O�W}aû�sʸ�~>�P�m9�S����^�7�ĶWs��g�;���)��;�moiG�X:�
�������ڪ�͍AXs �����m��
ŭ�rJ�I v�C��6�$�����4��_����FA�nyϠڻ/ճ�+�["��ߧv+����j�-h�L\YN�Q���r�i���Gm0eT>+^�-a���&�R� ���`�q���!�QBei�rj��c��� �j���[j!s�ޢ/F��g���k���a(��������<(:E�U�����1��薹���v-E9�K����5>^�&r�T���kSibu�+�ƻG~�c����e��o�-*�F�2;�Χ����>4�/W�&�A ĕ^����+��m͑�}��N��MV�<|�7�'��:���utzЂ���86	�@��~���(	���y����w�rH�N�H2� �0�%s�0;n�?��ϳ�\��Dv/��T��q��=I!����|˔B��ɥ��),h�]}�UF4B����H��ɘr�%;���4]J�9j����F�z���aY�O|�}���}�R�T����&�m.9V/!�����=(+{�P�FN�|�}�Nl�9�Er��\�����s`KG���W�ld���	�)̅K�j����&LC|P[HS�
��<ì��ϠE�s@b�-�ѷ@_��X��//��w�a<���^�6���<���2�����MD��d�0�K8x��GN�lr����:���F	 Q�ϠT-uT	c���� �q�i�^���z��d��k��
�[b�F}�9���e���ʾ;�(@̱�04��;��E#W,k��@�����]�0i�o?��s�L���Qg�p�@�UpBd��Jz/\�d���<�\����9q5O��ASR/�bz����.� �Ͼ�["�&���Ş,�j�}.����+��=��._{������NL	����g*�!�ަ���s�u�}7]%����Ν��ӹ�����yV~�,���{\�%{E`�m5^C�Y�U�5�5@�"o)�2�'�t����ф�$W���c�:I �5�)[c��R����#� �ȳ��DZ�+��"���׳����i+��1�%N�)�5K���N��f�0�}��U&T�N�߯LS��?��+cʰ�<�K���DRj��j���^��M��dT��C���:ֽ��%�E.td]�_{ݞ��E����O�0_�#�Z�V�;PeY�!"�3���a�lԇ�Uݩoc wy��u ���v%*&�&��E�c��_��ʭ��G���F�a���� ��1.a��hE`r�TsQ�
r�'q��X���WaQ�xԪ�B�� �蠁�B��vCk���"�f|��Vi͟,�����&��:���Y����;l�A���r�aSg��)�V��}���S�J\
�_�����ۙ����f���&y����'�����,���՚�^�+�<�*7�1M ʴ��VUQ�����ug��&��Kt�	q'EM�o�9PJn��6�C�;���9��B�$�.ǐ��G̱�g �Dqfj����]"�ǎ�o�P���iq(��W�'&�x�!j#�??��c��d��_L�9V���^��]i\(�e�+9�O�0�2��3n�*������e�%�Q�<��ɺϡ��IV�Lx�<��������u��{��H�^��Q.���}:A1�w;�)��}���iQ3m/r#��7���u�̌���s���gpo5����C�/�֜���v�t*<[<B�N���@����#Ⱦ������4�o&%yIZ/�1!9�9~7�$8j�e��>�T�?�tjJ6���t��$�:}���/[/�x�V���WN�'���r����H�V��S_�Q�F��nL�N�]Ѫ�Y�5�N(�U ��������i�����)4���8q�Xz�v��)���rbںku�aZ|�y��8�����hެa��B�NQ�A�������	�nȜ�c�^��Q�9 p�����������fB2�?^�߰��ڝ�C�~�'@�xd��0�n�"棖p�!�4ӡ���L#�q>�#���ƻ0*;�>����g�q <�Pȹ�!wN�� 	�����;szi�f�YХ���FC���hD���Y�R�cr�s�������f��v��V}s���K�L.冃���8.mι���Bt��uL}u�`�uhr$;�����lٌ�d[6 w�Eo3��D��vT�H)���\\��#T�����d��M��g����qO��,&���ﰟL�eP�vTj�8!N�vp_��m�m!BI� o�s-�Ɏ=^�CF�����H�a3!��[���/&�gf%�h,"�8]:P�|�m�n�'@��@�{�Ҳ��F��v�ӑ��*�f5�љ���?(Or{�f�7�S ��W�<����q�����mri$2X�S&R3i�H���Tg�5S��a�8T�{�G{2ic�	�|�ś$���Ƃ��tJ�+�TzG\�+,�?̷�n���Je[�[�3$w�d�$�7% u�|@Lǆ�R���}K7V[hu^���E��«#�ј⮲��4�)Y�S"l0��]dR�IB3���L���F�#��X;g{:t�0���Y�#]u�#�CKD2���0GS���>�ک�yv�馑2��4L�<e��E�jbcc��'�0�A�0 ���Hqm�Dk\���g:������4�K3��|���^�8Ɛ{<]<�P9��Mm)�{6���u*��P�8��lf��M���3S:U#1Xc���w�s��|� Z�>j�#�&�] ���w͝Ϻ���$��@;����K��^M%q*�P�bv�K�	u�U����R�N��r���ñ$^���d/�u�0��c;�4r����֧<������|�8|��@�7��*�����C���R+	�c0.8�O��gCC��%R�wV����U�o�01-�4��x�g��i��7�%,c��<���\r�cK<�:焱.Y"��@��|aɣ�	Ƽ(RJ�#�})+���B�vws��4]m	%p5{����dI|a;�m)n�i�����Tp��abą7�0b�C@���`�إ���О���D�4�P��&"L �E�߄`d���>ɮ
��%����/ %1�����wX
�KpX�CJ��%�WK�s��d����nW3V�nb��P����o��uc;O�%R��5|����/�[燋ۆƝ̲�#,6�Q�=_��贪��!L��.Ň_u�:{���E�#��7�0�qi=��Ⱦ�@"xq�P�O��N���,4���D�P��������{>�t�����Ⱦ>�i��u �<�e��\ҳ�(7�$a�d�t
[Aйߟ٨���JdR�	J�D(�	nݫަ%zr!����<UmͿ6�ڣ�exL�Q�B�U�#�U8��.4�k���܏V���I6&9$�WL�!��!���r��4����l���\c��'|x�V��>_ʵ����md�`| �{Բ��Jhus�	�<�̇�����g��W�<nB�I�7��^��y��7�~�S�q�ȄI����@H�[C�˅x�*����P�!C�2K��'w[��2�yIݴ��N���6{��W�A�g����cJ�ڟ@;��Ę�w�&4捋�o�m���l��_�$uXX(4@�4��tA:V
�3�޳yPܫ�L�S�t_!��M��}�[o{���7/b���ɱ�>��"��z&^��W�R*�҅������>vʐhg��A�zw�θV� &Ҹ�Mό�)7E�3�L�q^V���+B�U�v����:Fǩ��V>C��5���o׮YB��D��Y���(]�[j�6����5YfE*�G6v~3D�$l��ƾ��T�A#T�8��y�b�;����@`V�/Lc$�-��9?����q7��ҥg�z��\YN���N���V��d��G_�'ؔ��8��f��~4�Ia�$�
Q'Z�%	����[96Q����zD�-��� �����x��2T��X%p���b5(>H�f�� ��C<=���Zk��ɫ��9�ٛ�[i��^d�M��Zִ�ύE�S��I�uu64&�l�6D3��:�W�A�0q������m?x�(줃�W�uͰ��V�5�0�PX=��c���$?}���OI$�l-���ʴH,�
���lK�9���R�괳���&�QM��G\�\֏,?��i��۲2X����8j���,�P\�c�h�~ �a����uP����I�y��-E�`�w�Q�nR���|ک*�D������-��Z�ȓ�MW�i�%������g#��.	So+!{����,���6`s��=���%hm
�j0`��������\]��.l��ٲv�@a;�]r����e��Ԣt�Ῥ����e���ŨF����pmᚂ5��Y�_=}ؕu��6��B����hb��&���h���2��fCz9[�Z���=�1�D��Ĩ=�ꜞ�f:6�_�89w�vVY��=̀^s�w��[���@�%������~5y|m��,�ً��Lb<m���Y�wӆP�Y.]���v^����G���8��G�Y����`��D�.-��N������}�.9���h���W�a:;e�;���e����\L	<C+��c��'<�(��p;zv7��Vۿ�Ļ��Q�u!���YB\�"�)a2��͚%o��kP��}�0$��g3��?i��S>{���˩sA`����e����"-��t�����0�=��{�څ��0ϣY�چ/޷�

�U��ׇ�Eѵ��%�|�{^6d|(;�>�iY^��ιd��S��_D� �2����d�i�/�yh'�)�3I��f�'M۳�رH[B���%�?w���:��$�C��\kS��S��9X����ћ�&�/��U�q�#֫�BK�Sɔ��6�c#�Ј�e�iр�l��϶��3�����R�0g�}�|���5��*�7�$hU����eHe%�2z�	R-��-7��ȶ�i�T���	��b]��P�,?0y%)�d����$��F���6psVA�u�h*�]R��\f���� l���>��@�^�L�[�b�5!�xş9�	L�Q|Ҏ�Wr�!��<_%g�.�(�\�Bʌ��[�UA%}LM!*?�^���YV�l���Y��/�s�"��i�����_���pG�$����Bi�qJ�%�i��K�ҹN�<�6�~�[�?&�ࣲR�u�/m���{,���Rs��$��2��MB���_���!��v3&ʦ�0YX	O��ʙ��c��]R���.Ck�[���-Rr
���D��n���=X%����ՙؒ��G`���mb�&�:r�!�i���H���˳+S��(S��� l�Uv�2t���+�s��U*��A�4������LhA�h���s⢶������Q�v?�R����s]���� �gU^qP��W�B�ꚿ�oCI�rf�y j�'��x�ūTM*�t:Q5��B*��r*ġX��C�Ems���a�]�.c���,�ۣ1�e�C�>0D3�4Y�F� r�z�|b��gU���u'��&u�39�یU]Q��[h7 �_Q�|ϋ�_F�C����;c�&:p�(�d:�Ւt�_:f%M}3�9d���P�u����|���q{j*Q�z�Q�n"��u��L���Ւ%�� ������P��2���DhoW���:�F,/�4Z�+|�+��/P8@N0+��` �9��,�i��vI1z���8/D%�a��!bMB+��Z	�)�Ǟ��n���Op/	�G��,�N/��8���L�77V\�	�h���{����f�_���9����>�ET���53���'i�%��ʯ�$v�S^aWJ7g`t�\D��Z��w{nV��͐�(h$r|����O���V.f��Ȉc1�n7� q�YV,����{�B_��g��թ\����ܰ�;9)�TTXx��O�����5�E��v�N
Hg��� �q�eίU(�TMׁ�WI��e�4�	f�L�Jn��ӫ_�K�v��6�/���}8cE^tET��&R�A�^8�]��1.Z��4"$�ϊ�H��9�R�9`_����聙��:���*�^��F+�s���_&�I���r7�3�{��R=�����C��t��R����
���=˓`�Vd
k%o`C��r5�T�+>��kAukԔ��.X���%������_gO�;Tu9�n͈M�gM�pLsx��֌��c��o~�X_Q=j��&�!3�m<@r�F�~���n�֘�L��9��/~Yce�����ۑ1GP:غ��%R���v�q��w<�ʻK�Q�Y��t�u.�kaI���ZN����\ت0m�w�Vn�M�B�o+���5$*��+���{��,�K�4jp�CL���-rb���c�O�*/�8�?��ռ=*Ɵ�����*R3^� Q�b	6ZM5p�ѕ��C*���ؚL�ő���/���T<�58��W{ò���:��Mu���
@B��[����U$i�D�l�V�����3[{1U�X}���aW�E���K�2B0Q����8?
PDԒ�M�[WW�����ٔ�w ��k뀶Ws�ݛ'�D\���v�_���t.և?Z�F.�Ο�#���~�,��?����2.�}w�w2��<G�a���Y�t��ɢ�μmt�ݲ��� �O]w��\�i��t<jm�߽��@�፮#�3�\+����y���/� 0�������gB;�'�ܸ]�&��f򓺀׉�U	MJ����	$9��ӱ{������9�^v��W��a���M���M�>�_e�_�y��Hmd�W��k�d/��.�]���[|�bZ
�l�ؼkbG��.�\��[g�|�/<�~���γ
��I�[�a�v�U��0Ldg��/�'%�j���H�F��}�΋�[z�]Z�نn���=���ou.��������vG���p��WK��r�+���M[E���8D
��H��к��q�s������z	89;E,�)�N�>�P6/�F3�a
4���pϐ���Y���2{F�B�RmrB��{�jӝ٠�"�i��e�F4�&�R)�]����T�(�:a�,�qL��bAM��w�횞=u����,��د��s[��O[�7O�놕�*(S�U��)b��-rh��R�Ɇ�Й�x)1W6�o����(C+�Dg�5A����V�e��p�w�ن�65��oX#�i_�-%N}��t�Cg�CEz5O�Â���S+����*<��d)Κn$)�� #���|���g�Y����;�-�aA5;�]�d�B\b�	�59-��e�[Zq�;?D亿ǩW�CF�Ā"�����@&�^aq����ꍾ�d�;F�W�?o����x�ؾ����Z�6J���]\�yݣ��:Y������H��ޘ�����臬餪��%ԛTgPC'J|,�OT�;��Wc ��NI-Qr�#�(Yԙ��S�Bˇ�xT/tlZ�b�ހ\[�K�;Z�.�ͮ�߳)�j���V������jbU\�h*u������^ٮ�̾������>9�rN�z�h�8qtT��b�v�56�����8������΅��.U��~"SG�@��8��x�U�H�����M���&o�\t�{'4��\�����a���Ѝۙ����5X)��1?M�� ����/�N9M������M���s
>���:F[x��&k���5�s�J\k�Lw
Zcq���x��Q�xGe.�I���$�aZ�5�xj��������9����ǋhP�PI����*˚u�ϝ��A7$y#����렷o�]�/%�Th�׉k=��5�u���aA�ڎ>�T�CHB����Vٝ�3�~�N5G�C�o��N
Ⱥ~��5�l%����5��I0��@�{��E�q"*�Ci�Gk�C�I0�#�E������L.��O�8���=V_:PH{@���Gy{����і�Ƒ
4��P%l.L���O�[)�	��q	 �o���T	 x���z�P��^&>�puч3�!��\a����;��j���VX;�l*,��f�&$�\� }��skk9l?|��7W"��G�$�rx#u�d�Z���HNg�`
��Ӱ������˪�0��@�j3߼$�Ø0Xp	�aV����qkK�N[�6v��W����������#����'m�"�a�h�@&��po4�Le\�)��[�+��۔�2�#F)yv|冴{A/h��mꎂR&��Р/��X�W�[�X(�ͫQfH�V�_K'����ߜ���5l	����� Z�>DT��雜D�AF�mP�Đ�)�M ���1�0�Rx覹�9^L�/-�F�
P�Vt������t����t���p����h��M^��j/���w�Es�����!����[��V��Q(���IH1%'_ιY�4����m��瓜��G`��*������9��M/�dT%�Ø�Ԋ��_U|�v���I����\��@�@�
���9�<]m/6SGdy��z�\e��e�BZ�G�-�#��DR"�9���x�%�nԭ-ʫ���~S�T�^�e���0{S�p�3Q
�h����}���C� �\LO��y�J;KLT*?vk$��LW���ט�{����|[��w��q0�����x�F(�T`�.�4�:���l���黋k''�ڐ�b)�!�t�U��#A��FH�ٲ���Z�T�M�\����WH���d���3�Q��=ׁ�Ụ:�� N��~��s]�B	&ʃ����)N�N�7�䌪7NI�Y�G�?�Y��wS��Lg:2{�i����f��t������;؅�$S��Z^�Y�5�;���x�E��B�泄H;	Ac�JD*��ͤ��焨�v��mY�~�{��zU��#6���:���Qг��v]�L�}�uC�����9<+
��zj��Y�`�� M�6�j!�GȁcF�x�FU���!���w�t �#��y�O�Gg8O�V͋(w=���v_���n�bΡl����LD���ⴿ/:�e
WV	3��<?�ÎM���p�qT/���m�L����;5z�a,AK�q��8�Y��v�^�N�N_M\�� �%��U3���j�S����DQ�O>%��+�)���چU�r=[-FB�/��@�}F�k�?̙�Z�x3���6�vOenm[�@	�y��!`��|��k_i�/,Ts�
=��r~�+P�}��I��A�����)�!��4�rR5��edf{]w��@]鰬ΉCf�h��&c8K�p;��F/+nG(47�K�G�m(���1�Gv�Rd��ʂ3oC؊�e���$�爩SA����ۙ�G�s�~�������S&3j�l�%n$���X���̻e��t%jN�<�������*j��Ha.�*��h�~��T{U�Yyg�@�J,�/� ��jÆj��flg�
��D�����b^
�a�Ͼg^Rvmu�C>'�k~��e����HHXFcH(�~���K�V:~����n��U��dC�yH�Pz�I@fk���jl��EU%3�z���֑�^�hld�j]���Rc$�ɖvL��?���8C��T��� ��I���T���߬��%q~*E�<���ֻ�@f?�[���d�HFz���2ߕQk_�����_��ɣ�2?�ԓ:�.��}��l,U�1�%(S��u���UC>����q�h��T�	߁�l�#�*�Trڸz��z/�tglPw,�e�΀.p�����~9:�VDXt�WURm�Y��R�t�~�ߓ�p���pG�8�T�F�^�-�����Pݏ��^[�������SnF�Sv4j�����Z�}�Q��af��� ���=�tsgV��Wj�˟"!���|okx��c<��%��'/�H���o����Qɼ��!�t�B�鮸���h�~�&�|˰)���ž���I�޵{˫�����O����[d�	���}U�C��Ay�(�*��<��s�
E���+�.qg���ԑ�gpOM7���ь!�z��i����q��׭��Hd�%�]�8��d�8���ct֯�t�aykx,Aٶ�rm�x<�&�X�͈Ư�!�Iahm��"����#[��ݝ���I�Yk��G¹�N
�d�W?�cA���� �h4��n���_��3��BlWL�o�����7GQ"��d�f��zR�ڻ�D�C�0���%���WR,�c��眎gS��lV�DBm-UsN[��7���4��Y5����h�>�ǻJY	N��_�}��*y0滁|T�IWJ)�����Z&�M�f̉�̈���l��HH��gPf�px ��x'�L��sc����}#���N�Hb��`Y�����8=�u`a�/�,^���_G�k�r0 �L(	�9�����ٙ0�?V2��~���.�MΑ����պG_��]}d�A�m+s�}y���dM�v��:1��(!��s����Ly�x��{���kZ��vMMT ��_����'��J��I�z��B��%Î���!E_�]-���D4�P��n	�ŏ��'2$:�C� �g�J.o9�^|+7O��WW ��ײ~�^䰧Q���n�CGN<���s