��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	��E���Zګ>�(s_�
u��>���<Vx��˜6b� ��<�T�m�I�
z�/N��4#Fq��5b��͜wἦ�xhaa�PR�,l�+g�L��$���Rm~B�qg�o�
p1�pC�`D*"�H;��7��:`����=nU�nb����cZi':��}�A���'^�8Q��hz�`��*`�GO����}W�| ��N����jw}���h���;���ǚ��0���:���X������`�[���J��%L��m�
��V�e��O����)%�x����JݭW���<p�[���wԋ�r[y���ȩ�zd��!ш�?@��ƙ�V�d�U9�=φG��Ja�)
*�/Ps�0+��z�ĥ�k8
X��H�ws���QC� ���KK����t��Km�?Ǝ���*�QQ�/��d��+�x�O�H�#��4p�v����4�9�'�aPzS����p�����$(���u�����+)|���S���OT���^">�I�S��t��i���ǌ_u�F��=|�`����n�u�h*��DN��R`�;}!OHC�~~�N��%Nid;����2b��6���|VG�8O�F��s���
`|ݐ�@�'Ѽ��=����_\���8/@i�f�^/��)��B�#��ʱ�B�-�4��y��&y.)�_�jd�I��F�fx(��˖�g?��d��@A����_{���6���0�=(?�p���1�<�.�# �/5��F�tr~ տhyo�x�s�C�e��0��@��9e��u-g��A�ށkA32��=$�kb31N�΍х��;�k3��7E �:��Nɐf)�����_Q%�\է$��~�`�7�=&�fĨ�â��_���,��4Qq����{~L
�]�;���u�6J�N<�&�)1�!Ô���e��+ݕ���B0�m�7)�Ke��&䔐��8dI���(���:h��k��s�bM?���!��#�`��Ĕ4� [���z[ݧ:g�l�Fۭ�i5a�v�!0��W�Sf�`,X�3=c
�Wg�_���Q��Rw���j%Ҳ`����%0 �U��^�M�d��:VHT8��;E��9�wnȌk�;1����=(B�<}�h��ʪ���O�!�a2I�D+l*eD�ġX���vÃ���Hؐ����s��0Z�8�.��yd ��&R��3=�F��U[������s1S5DBC���˕0�~��V)�� ���o�Q<N�P�$�"�����Mx(�y����
 �,��J�2hbaY0��l*�����۟�*3ތ�]����N"�dHPŇ�p��u�r�F@2ؚ[(3
ӟ^�+ɜy?����G1�P������>�����p��   ��I�3id�#"���������<�[�b`��x|zV���D�����k��M(P��mfgG�@��U����N�}��{2f�?�e���8X@����d�A�����}0��$ʃ�W����A�֕U��+�WPE?{�.Ģ�*� e��{(��m%����=x>�a�g�[����B_�-��Q?*�kU;�� �c2�$ѐ�q�A����T+�%�*���`D�Țq, n�%Y���7�-M���A�*��I�@�Ke�Y�.d��-�
�������O�Q��J����%�|����8_�5��į���}��E�Ժ�«�4r�i�..^�>��M{୤.B���}��	�*�9y� `��6�M.s�5���܌B�,C�(.�xi�_�7�8*��۳�1m�U��K�G�Օ���B� )��|�E=���	�W��cp$�-�5Iɺ�8��B�Jut7'�.��M�B�����Ͳ`�U,B�ő��5��D�Wi���!GOɥ��4���UҼ�6J;��63��|�[s��Qz`� ;L|����'xC�nʘ�T�OOQ?޿̻9��;��,�!%�D��KAv�Z�؆
@�{^�j�JyJ0pqxK?	�}��*TpN�6�\��sfdRx�{#��0'����Տ�5�,/���{��f��N2��q�0~XKk�L�K��n�t�����*0M����bblkZ�}5����Il�ԟ�
0����"kN:��<�?��8
��]�h#�?tǿ��	���ҍ̥����q���㮽��ou�O���&�Ή��/{t��6z$a
����ޣ�"�y�Q6 �TVĢY�el	��ke�}�z���+�����~�ݸ�`e�fZ�g�qt`Ms��o�r:c�o^���,�'�˥؄�"�rG;��p͙���Bi�	;�E�qA�<M�Q^,�$c�@��/��+�i܋��!ه4�Fe��]�?\Z�4c]�kS���L�qY���[z`�`����+�m`^�@�x�(�g/q�}<g�CN�#m�d�HI l򃈱�o�<�@j�8b,���lS�L�F��=&x�蜽���gu��0f���x?I�����\�7D�sf��૞�>bT�\�l>}M�n�v��'�^�� �R���-2C�iu�����0�8�c���)T��ݱ)�?N5W���(f\�m���ómVhť��{�]�,x��q�S� �!��xd7���@v8��)��"�]^�ԞD8a���(��ʰ�A�^�n���N�v��r�j���x�+V\��	����U$��g��ONMFk��c�Q��~O���>y��[�RƢbU����Y����'��Pc9�h�Pʯ��ʹO������1���L6,�~(	8���52>��j jx_V�a��s�h�����:#'M��?�ͯ��(�e�^�: H�E�a���c�,��W��I?�Vlw�R!��
�$?�Y��P{�+=D�o�uɾo@(0�c��vEJY�����n���(2U��e25/|�O�F���zE&B�
*"�P���\��ӡ.�ρn@^�Jb�� 9��0�t�Ta[�҄����U�֥'t#������e�"���۹s��4�����ݻo��L�Ɲ,q�@�F�%�K����*H��9�B�<ǚ���u�,ӝ�q�
�7��q�w���fkѢ��h�X�k�m�IW�:�uN	���%��\�?�Arw�J�����pD�2d�|�x=`�U��HA�:�g��Q~�	�wGkӄ@u��{%7[�W�����;�j�pl7��*��BӋ�QH~L;�_���^��(�G����y��Sma�� J,��2$�7%��/�-�9�`�("I���� Y�n�I�+8��>v|KM����֎&���i�zq7r�������D��R�������LxN�w�Y�&\U%&��D�l����Bz҆�jo_P����Z�!G��d���5�K¨��Q�˘�_��&��z��~D��5��ɓ��<*�2<u�7*A���Y5Xl��j�?Uy)���/pe��#6|rıho��G4�
M8�x���Y4 K͝n�n7���%X�II���X[��	��jk�)�b\ׂ���!#L}c�[
� O�3xQ�&.u�)��
J�U���%�~n^���^���\�D����n+0��j ��À�0��r"�$^"#{����":e�_q��`��%(Q�� 7g�S�( S�J>�t̚rc�&�ݞ6��
��y ��	�=�{�h��1��o	X��A���*!H�F�͐��Z����aయ��T�xӟ~���`�b��~���@U��v��e��V�l<X��=�>C�/=��$0`0`��:��N]Q���%��[�����0\�f�Z-K�O01�Cս�ը���̩�&q���2;�u���(YP�t9��L(eL��A�;���6Z�9X���;�U��F$������{��}=~�24HÛJ��ݖL��'&�a��
�&򓾐�]½����X
�-D��$�נ�g���������ݭ���ji�.��#�E3�v"���Ë���K��ں�<�@7er�o�"�p����gI�d������6������gq�u���]%L���W^(�Wj�M�*���y4rm| �T#�
��6�d�h�}��gQY��������bK��ڐ��B�@D��y�nv��1ˍ����U���r�2q$�N}��3n����jv����p�	I��T�i����E�
��)�]��e�<Uv���D�鯩_�X�ǰ)OĨ߃r��'K�5��>�rub%&��E��Q��| Զ�?Nw��_M�D4��P����`�B��Pxi����`�_/��
�	c8��0$��L�S�p�~b��fh]/�b������Ky����gբ�@�%Aʹ��AQ}�;��z<Xt.�$���I�I�?���%�"�{�⨌�=�vЄw�u/�q����ր��5O�<�׭�ݱ��D�CZ*1ƿ��Z���F�J�;P�cAC@�:�j��G�X_7�(��a�&3nE���Laָ`PO2�@�
����e�����+>�l��\f���J�(LE�$�ƳHF�������Rfl{0���Y���a��탌���3ܔ�E�5�_I��C?��A�?r�zi�;��C@%(�}��Q��y�k��7�Z�f�����%�섂NF�!���~�O�x��M����)"�-���F�!�ɩH��W��Чݐ�TPE;k�Y7t$��3����\cgPm�5���W�uK��5.���s�E܈>W&��]����ub��4A
[�/4�+R�.��{���_Dɒrz�"���;/��k)oj^�[�� @:�~N��p��7�>��a�c(���e���� ��[豄d�F��������L�Im�\ـ�> ���&�\W����?��la$e8�>m��M�˜��Be<H��ϧ�K?7�R�;�]����F�}5��&ך��3��I�l���^��1�' ͚h���2�Hb���W�����CCxT8mP۹F*����:Z�x���ڣ���FU	Ʋ%�c��	�j1����ӑ�:��m6<� iS���n���ӚU�&j�xo��R��@�d�id4�2h�����U��kp��IZ�J-��&������yq̷H7�]1�|d m�-���G�g�rcQ	T��}iB�o1>�K�b���RK�XN������VڤN�ZnHս���.E��N�}`��7�+N�/D�`3��4L���]�Ӓ��������4�xz��Qw��nL�>��Bn���,�l�mpn\��,�Dnf|�*����<�a"0�6Ǝ�؆��6N2Ô�
� ��;2O�5.�8�����S�b~��*������Ya��z��~Z��n5�<���r�1��ꍝ���(��ߵ����P|G��:�8�֟t�����ǫ�fʄ��,ֈޑ���sU����۪!I�\-ߎ2g�k��`�-���j�DuO49��m�5��$v��,��mY��CC�����&vz����� ��K���t�8m,�WT���'�b��+S�q�%O�y�`��L�I�w�?O�q���ۥ�Tk����%B��i�Kc�2��q!�
F[d���g�cZ`�7^Q���q���w{^c�k�8�����11����y0�*ʙ�X�؊���k�5(W���/D��0{�?�ȕ�����Vc�ڢ�9��mm��ک�zf��ΗX�Z�7��աB[Z/(j`xYY��ۮ����U�5c�4���<����:u+��{���#x�|��K����?��t��6��G����|�%�])��³�p�P埬�q1ļ��Ͻy���>��ƙ�պ(�niqURV�vw�p�dY7}�r�AAY��c詅�C���3����#��n&�V�	q���P�Ȗ��)3�q�XB�H�iZؖ�-�HD-k�fxѧ[� (wb�6�l9�~��	q/�2\�n����.M�������GРP��-ܥ5���&V�����`'ۘ�`>=A����>��c�����5�����3�dZ��P�n��f�)?C7�/����?nljTYx��ۯ����iCQ��@�x�e�O�T2�C��_>�_To�QZ�C� �c�.�U�"dY@ԣ��m�r�C�m)T��~
ë���9�nJ�ĕ��?}D���'�_�B�.V�Vm�_S �+nB'��ٶ@�|6�G�6��5h�(��CqEI�li1ѕET5Ѳٻ������F��~�ږ娉L�?��阧d1_Q����a�È���u�s�*n��sY`�E���L:9�e��D����e����YU[z�I�נk�Ӗj��'t\[�V���$n���s���r��o�����L�z�95��~r��0�v�y_���G�c-���脩�l�ω�6�m�a�έ5��v�Lq�S�
B�7�����.�
t��]���$�'r]���#���U�(�׽ �D�~7��<��B@������\=2iX?��QM��M��.�rq��1>�mr`�d�՗T����l�4���X#��#��x��X�Iפ�慕K���.h��`#����L�����e�H�*�5ݨ��I4��K�Al��m����os&~K����5d�E?�d���`Y&
��}C��*�+ �Vw�j/#��js�m�`2$3*���/��_<7ң�:obT���u���$H�÷���X]7��&i�@������l�S�y26��ꪅ`����~���ۺ���7�3/�͠�
h��KK<ʾ�����ۨ�9�-�8��SP��*�V��t�ؓ��`��:&}^����1"B�?�L4ө��ߦm��Ӑ�)�Gu��aY/�f����^��J#t��M�	(MY�\�	��"�N*�\�a��?�w�a)y�wG�	4XDnQxp�o�Yu�<��9߈�3ߏ&3%�~�땾�[��{�?ܝ����	���������Qf�k�Z�7T��u1�s�%��v�js����.?���3�8%���4-NEG�~BF�e��+�k��-w�ܜ�l���N�?U����Э�d�	8O(�������(�}�0��"�pF�N�v�A�9�������5.��̖��L%ԫ�'ۯ�������'����Z���#�o�ݓT���祮�ݰL�i��S�c#�q��+��L�V��TUw/�<���~��d�a!u�&�(��:f�*�w�U���W0z�/��;͜3��N?�`>�FRl>a���	�/v�ʮ�ٺt���>�}��}�x�u)�
	�c��N5"	!�4�Ku|%����d�;1��\U�X��]i���a��?�ox�S>����VL�Ps�B)��B�t��2���V�
(�����5M�r��X�Ө�4����W/�p�:�W�u��H��(y�t�R!	(�=n�W�u�g�*l#�Ҵ"�[ɉ�<����6�(h�}��,)i�{n�z��{��H���eⳡ��Ųu;�	;��;@�(�P��ɳ���{�������&1��WZ���)�5�GC�{�bd�H��_�wۦ�+�>ޗ�C	y��v�y�f}�.1��l�|�,�GC|�Ql�OrY��-�2b^�m�(�)��ӯT���8tN��_y��!Z��S�� �Z)�]�y���<��0V�Lە)��}DU8g��=�	P��XO�.�����X��x��j]�}��W�|��>-��b��ެ#;�6$���)�V������#�7�oOIM&zl���jz��;���T�fJ����_��_�y�`2�3��(��'#+ӷ�j��
a�Tq�@Ӓ���M�E1Ϫ��B��[$�F�^Z�CV��$l�K���s������P{��ļ=�X*X��1�f��]�����H�WS��꺓�1��F�hK������ɔ����o�}iҗ�0��P�RE�N�%N"��J<��\�	����A}�Ȁ�S��!�YN�g�(�0�T[��{&!��}��v丒���n[8�{��Xba���
jC�K$��3Vl�X8�n�vj�6����_����N9w
�>mG�ʹ��yN��i�)�˕\L�.��eauo��.WI�ϲ��r͔l��
]�
�8�X�Q���O?۾N�Z��&(􅧌[�s�yr���� Ī�>Z9&�ѡ�w"i���8]&���xBя�jPO�Th�}$�,
���&ݟ�}�b��	���R��ȴ:(�t{�б�)=�!�<ږ���%*�f�$�:Ș�@��)_�e-<�e�*��LH�Hm��S#�oyIw�䃤W�se��Z���a<���ߵǊyZ��TzT~{e�HsCF"�@X�K�X�4Q�Qs���;S��ݍ�mh���Sw���\�n�؅Ix��^.w���������{�cscJ�@�~w�_}���O�(VI�(JK�1%y$�2;���7���Y��j��۶��x
L�ߣָ��x�:('�#j)��)z�Q3��
q�e1u~���B?�����ޔh{�K3Hl棹6�q��[�-�`zRS2d)�\�c6J�fD\� ^��7&�)f>�cnw���9=j��9��4���*ÀL��3���̴t�&P��X��+*$��EK$�%��^�U�N�{�r��)Y�E�c��ݗ¦a�un�q:��Ty���\��z�v�񌸥����7�>I���JNo9�M)�N�m�[��i�]'q��n�������6�{�|}'�*N>�O��}�8�V
n�텩�?��Б��k��/�+�	�5��s�����:ą����jx���V���jT-�~�����
n��NwEF&�ԝ鼓���u/ԣ5�B��:�C��Ǽ��>,���b����=P*k���q�Dp*y��B*_���5��ڮ�X�t	XOR>3G��A��f�Z�]��/D�ɷ"֟�c^p4~z{�*̸������[j�f�X@�Mw�}RV�h��<ҝh�e��m���~ԙ���_n�������jvd���7�&�=9A��k��\1����w����e�.�Pe�TL���֜Z��`\�f�\Q�Q\�}Ա�p" ޚPZg\ �r�c��)�(�F4�����Q����^�ig��HSnL�����6��:�M��P.���i�e
�5�e���P�h�.�;��v�7n�mL�@O΂����2���K�@!D�P� ���x?����g��&��;��p������E����ɩP�����;��g�t�9k�Y�A/��f�B:�X���-�������t!{�2���ZW$Q���o,H�.�D�Jp�l;�h����Zb��&�]�)�ۍ)i��@�2�1�IF�\�e��`�}���GЎDbā՞)�6�^Z�o����r$X�:�/�b���h�� ����c��r��k2��!�y�$L��S�崿 �Xȴ=ac�5�_�v�XS�T�����JT��)>m?h pm������a�� BU�Q-��,����?A�l�z/�Z�x\0WoH1�c�K���sO�����8���.8��	�6��jI�9�d��$��;u�hK��7������A�sgy�L���G�ip,���N/�{O�˿F�w��;��ǟ��Ŷ]�7���wMP�O`&/�=p.e�����J8\5�;��Ԥ[F�I��a4�"��=���l��H��O-�������ʃH���H�m�N����/�Q�����/crJ3s�t0��}�J���i⦝��7ɩ]X{��+N3J�'c�UI�+'�L���j�϶Wmˍ�����i�X�_�j���^��_�N*ֻX5Q�6����!��5�$�#j�s-�X��~�IZ�T6��ˁ��LY:�zԃ��j[�'3I���P~n��f��{j\h�����Ut�p��_q	� ۔���M��~��6�t��
�F%�&L���/x�c�c+[����{�3 ���<�=�ܚ�J5�4�E�u��2$�eA�A���9a�ĝ��Z�p׶���Z��7	�W֝�"�D���p���:Z�֓����U�nN�BA�gQS}A�b�(�j��/�*�7��&�)�����(�|��Θw22���*����?�q3�Г4W��>��3nt���_m>)�T�8��#��&�}Mef������3Kmi]w�E�Pn$f���|��E�Q��C�`,�%��f���K$�*�,.
5C)Lޞ�vИי�v�����\�z]^�~ֶKIo'rzi��_��GJ�/U付p3�*�:(6_</�������o�T[���5���{Z��<[��\ <�n��E�R����}�`��Ju/?ح��S�v*���!�R\j��!l�q�(�2�E�S
�S�9�IA�����q�� <7��F�b��e	��ٓ��]
���xT�D�������d�����rҬD'U�+z�a.���& �JR~mN��������4�^~㿣[tn�����*d��'`_+�mbFys %^�[�Z/X@���~���T�Q����duUXZ�٠aa�v�u��y���	z8�b-P6fZW֎��2�qZ�}���ZA,��|V>]�" �17煥PF}��~fb�J����O�|��@Īi�8����F�=fR�ћ���# �c���W�-���^�$'[��;��W�[�!��8���1���vB�B+��䚅Tx���+�g!� "�f�~&�L J#iI[�H�ow~z�cΪt>��&j�5V�[�)X�j���䖣�9ެ�"-B���Y҃�&�WZQd̍3.�(7����5��J��eHRT��F 2�ȃ0)i�a��K��O�(|�]�h5�Ff�H�<a�_�_�f+j��a��X��@���3+t�%����* �+]�{�Z~b&L�!vq���B^��;x��p��<�	���>�"��s����d+�OCJ������[G�j�.�`w��c��"��]r=�X���#�o#;���:��v(�1>!@����l<�)|=xG��CW�0ZC�0·�Bތט*v��=7�i��ؗ�R�����FFvjh�m���֦|Е�s�U������mh�����T���$	�å���Vȧ�*\��^#i5W��;:થ�(�`2���yV���*gN��\k2u��xW*'����f� /�Y�G妿!Q�g<��E��YP�m8Yly`s�4۱��l��=f_C�H�ū-��W�Eְ}�8X(;���a`���Y��B)��/ p��O�?Ç�e��U>����n�s��?$���wM���<n6tBu�g9����X~ʒ���`�7Ƈir;4������?�I����b$�h�^@��0�u)�O�w�Z9��L���3ї�ղ^�hsH�3�^w�kx"��w��G5rj=,K��DL�Ѿcr�%1mK�_=�&�Mk��[_5�/�<����|�U�X�!DE[{$̸ܤ<$���m2���VO��X�O��E���4��L�,��
f�����I2�"��[Y�(/�X�%*�SӔ�P��q�d��hX���9�8�R,��N~4F.�><K�Yr�n�U�3֜�t�9󕼲Q�
��nY�=:�ib��%��B�Z���!I>�����U��d��V�;r�Xd&�qB�� �	1��<�����*�� ��{O����R��qx �[��H�|�<k��ן��|Y4���ͧ�w,��I�<
^����� �L+*��l=;pB�Ё$��T�Ll����c��!S��}o����LYN}��EWѯ��]��\����S������������|S�����h%RX�2B��;$6�l�vn��O���~�wE�6�]��#�{)�����)u�uZ�$����῍�����,��lB(����)�B�����m �o���
4�6T�	�vGE�� ���@��c]�rFb��K#h��/�B��ۂ����\���O/���nM���`;��	;�$G�x�F�q�y��6�,YA�O.��m��jX� =䪧  m��u
����Q�V�H/İy�Qa��ȓ=���f���.�	��}3���Խ��ؐ��7Y5�#�k�>�b��w�j���c0�X�� c<˼3Ƴ�����F�}�9����,:[-�
c�K����T����{2�AK�H�q���x�j�KC
�%�1���(X�I�i?֬�p33���V!���}�Wn�I��F˩��`�j8'&5TnG�\î�!�A��6���(���i^^�2a��� �ƙ��y¶���*���q��l-���,bJͶ�ڨ5.�{�4��q�il�00�� �v9N���]*ߍ~��<U{�`� uX���\���O1�̫*�B�m/��l �+����אL��r,c�����RvF�z���)��Cn�qw����'dE�41�W�R�lz�<�Ѣ:yx]#��]F�U5�*�*G*n��0*1��t
.��\�-�~>=�(B��ϗh�3  F�{3����򄵱��L�p�)#ꄱ	������=b�D��]��s�v�f:�0�+���R}�O�8�$�d����&'��bї�έcj��G�&v���3�@�)�Yw�;!�t��rj�!�8�ЦP���o�U�n���G}�O��8?IZk�ؼ�sƙ�S!/
��T�L��)�_��;�y�����l�����[9����6]&jǻ:>M?9˥��^�
�$���BBQ新��K�f`,���}�ex�
3;��j6�m���q�t����s�y?���{�[ʒS�v�-įQ���	X/�0���3���2L$I6j�D���d��h��=_�zܓ��[6"�i��)�>Ze1�Q)����7V�	M�JJ &wk%��h&=1�X��#�\�@���H��k�ɡ�^e���_�іy��JM�і����
-�v?/,g�_���iΌ��V�ic|HԻ�j9�Z*��ilE�s�'TW�B�!�q�h�P(g���2e���镹��8f�¨<�Ha3*G�Z�E#��h�����* ���h$�gq�R��]`×w�� z_��@p�,d����Be
d8sIll������|���b$i ����e�z��r�I��j����g>k'�h����E�DὀљV?���1_��m|0*��Ũt�iS�,��c��^8�Jj�>.6���W��$��q�P9tv �&��c(�a`�!�}mg,�U��H��*����!��'T�#�gc�LD���Ӎ,ţqK*�����IJ�y# �6 �'�2ErQ`�
�3���O��"��O\c<����e��(Jo �����q��|$��zc2�T3!�<][�z Mԣ����<�w�
,l0���/�9D��(M�c\w*�T�ƛ����Z�vC��GdJ3oiiLd���P2%�\��y�k��,��n�B��8X�s<+�m*L���Lh_�� �����T���)SuE��	�<�Q$�II~bB���"�Շ�i~�מy:8��a,���v�uw�)���m��� ��5g?7I�p�c���rZ��T��<��JYs�k����d<��Q<׋�1Ua�h�I����*��E�/��	��Ա�j��O,��������3��<*Zv�\��bW ���4�����R��0�p�?Ѧ� VgSX�+"~U-�b�g_jZ����]yMg�KƉ����d�tD� �mp�{=1��jLeA7j6P���'C~�0}i;&޼��Cw���b���9$SIz^a� I�.`��[�^)���z���n��J������z�$}N1��y4�g���ޖ#�R�n_Ok���$L��gkʍ�X��z�����R�e��p �x�=#坠m߫u�i�n�m!���v㗻�V��QUF���ր�G��?�E��p븽+)@Ȗg�1��2!�(��˽�Sza�/NI�ٖk����^��Y���Q�@�Cx2Cf�@!y������ ����FZ���[�+v,���z��eP���d�o��Yq��^x��A\���x��4������u\��?!�HZ��ts�{T`S��c6Ŏ�Z3+�1r�e�d�?�I+����p��לܫ'���m������1GPB_������ηd�І�qESŗMS���c��9�J��d�RS���CQ8����K(��?�b��0�|h�7t��	'�F]X>D�5ykс�K�K�߻�I�it��C6�q�6�2��&�6�?_��vņ��!,u��s/Fo����֢>/Z�>�9o����屔�~c�M�����|�iy���-0���"U@��������5!& ��n�
U;��i��Haf*79яQ+O�&r50�:�m��5h��x��V�����zM3�B�!NS��ӗ�F�}<e��-	�?W���$�d�/g��z���I��Fr���:9��_�*�nU�m�bCs\2l�s�i��0z9�.hA>6O��/�`�Bw
V���Z�-�-��HB%�-����c��IY�%M�]ޔ��Wč]�4NQ�������8)�>�LV-^�t	:�P��jا|2ŷ�M�T�zW���Do�� >BM5ST��0U�e������9	��q�&�I�[���k����^&�H�|;�S~���*�fӳ�9j8��vݐx~#:�v��5�`�c�<��$]eS��Ά$F��{ɾ��F�-�B�:x�e'p�H!�$�8g�B;9�Ft�-��&Mz��P�x���Svok�b���WQT����8�+�:��
*Fm��F�R�u91};�X�Lk|��7a�d�>��)w�����51-��3���U9r#�{=rm|_��\iu&_&�՗3�"�2!���������?2G� �H���r ������
ò�~�)�_��)�fЮ��o�:��W�,15N�^���U�����������g�e��T?�"�)���������K's�4V�m����X�I����=���ae�sH��i �d1�K�ǹ��&�(�Î�d�ffs�Xx�ό�-ٽX�Wծю��PBp��Z��e���Z��"HXy^q���t3�Q�����ƴz߿�q���3~�
欺(�1�~��2�%���h����{�y�*Z�.g�����o�%�-�	x���dW�X)pʝ�}�Df�w`�2D�%��%���t;�B��zg�V�Jt�'�AZ�Y�g.,�N�mh���st��bz�Ai
�K���fgdj-[�w/)������a�l�^�״�`�=��Y� �z�����j-���_�g`W���#W�E�'A���v�E��BO(&�{���H�l$�jy����ï��_���	�كo9FE�JRI榐^�o���e����l��/ι�k:������9��4���03'���\ݓ�srJ����'cp��KbE�}_�:𒬀�@��s�i=U��8��
cܛ5]���w�?�)4f^3F��X�13CD `X Q�Sn��%�yf�8}{�{ꄉ:M�A���&Zn^��0�C��Ӥ�e<*M��|����l��O�*�v��Ù�!��Q�$�^�2j�j��ԗ���<$���<z(C�A���d���z_�0Eத�^P����]��W�[i�����eT�n�
_-�<I{�"n�߾��ׅ�]0��`q�g/�徏��n�6ػ���fd��*��n����}����^舴+S <C��2��B��,9)&KV~w�c<�c������V�Vu+�a.�:��G��=���F_x���Z�t
A����+\Gg����EG4b5_��8��{�Z4��0ɓk�&���(^�MaPE&;�H�+*�-mz�@00vQ8I�u0;�H�R6.PZ6<�cT�_���%�������:UF�`x�(*AI$F��݈�#k��ƈ����<Tu�_��jF�E�цĎ|Yy��VI����U���OB�� ]�!�3@6aZ�	o��]le>Z����ǩAM��nMQ�kG:N"@j�t�o[{CS��	�>m�c}RDS��tޭ��p����|]���7����q�m�)R1�y�ΨuۉB4���g��d��ܗ3��OM��_�?�`��I�A�	�v݇䗋p4P/b���t���,�d��El?�,��1�����YP}Е�
�����z;��34�_�6�c9�u�8"��<����B�0,�1?rl�R���4J�=@�~K�W�rNb4tt���vu�u�왜�����U�b.�M�/w�����tY�%m���>�Z�xm�o�Q�U���ܖ��6�bqI��Y#.�f7���5��?p���!�E�F3>L{�k��!����T�p�ʿx��@�r8���ϓ�\��S�\F����Al���-��B���� ��';��p�Y��6��L�Q]eW��iB3s¸�����߫4<L*5[k�Z�_p��TXvZ}�����p�S/g�h^�e/�����g�kOv����	����/����'�We0'4%��pR#�`� ��������й��KUg��c�{��P��K�q���j~���)���}���yۤ	yC�5�n�7�,1p��B<����C"���*6���j�&Hʅ돇,�����y�1{��T�k�VB7R w;�b�TeW@�F}fr�rxp�Nec%��m��<n+�.�잲q_�`��R��s�o�� �m܋�T��V[[�h��&��\���򓉀Gi�a�/�/ن'��ۏ���::Ҍ9��ۜ/?�jo�Ze}�2�F0s�X%������\e#	�"2?0t�<���f���a�s�N�	���NER �#yߌ �Z��4�
��'R�5��h�"ҳ���T�q5Ӑ� ⚧g���R�h
7p�9�A5�x!�C��N�lΩ"ݙ��D&u	��9,|y���F�f�Jb=͙�є+�f��j�ť?��|��m5�j�lDWY# �!RN{ �̦��B[��蓯����{���ܶ@嫽B%F�u>k�@�"���mY�d�L�|�-�$�ث�Q�F�hhA�>)���b7�����m�3�>f����8�8�У���m�����"�%S�os#<c������1Ι)p3����F��B]@�u^fݸbئ���}��&�%5��{�=�����:`Q�5�4_᪽A�]p�s2�y���\�41V�q���RC�q�ʗ�٣M�C����9c �.~����NɎ�nx�4�ͭ)[����Y�nһ��()��Z���؅��l�������˄��1v�85� 'R�o��`�Gu������JK��&A'�Ǟz�",  ���`������H�w�t��$Qw�$k,a��qʿ���x�_�y6k.Uir��)g��>F��Ϙu�
?Б�������;e<P��#�h*>�)�Ǩ<Ye]���5�#6kڧ�j��C<Aa)n}{X�`�c��a8��-\�����4�&��}��؆��'db|9�1���2?�j������3��ZOEY��%���h�Â���F�>�PF�n�X���?��wh� �-��u�o��]\'�x�~����5��xi�F�:)
��]�,�����Ď�3����NN��X�.[d_G�}̴Er.)&~Qy��v�E�C�Ē���G�bk-�`���V���k�XG:�q
�V�\kU��`�P䤿����L	�Hv$��#�	+�(�Q�:}u�v��%�-S�۠(\�OR$*!���੼�hw{�a�d�N#Y���O�F����OO��k�ZA���\Sy�!W��Q{���X�&!�+5�q,�T�೙��A�ivwП�A�
���p�
_��{�����;Ȯ{�Y]�������vyP�7N��c�p�t�+ �R�q�%�8��CC���(J���������}��}�-�+'�mV+��w_��e4=��L����	��\Hs$�P[F*E;�^�}��љ��"�Ijű#��M54XćM�0�$�mА�D����ǅ���e�A��[�h������V<[d�%m�y3?Ǡ1�$�'��?�h#���#մ�G*��"��wZi�Y�@�=��$e��	۽è�n��>ďHdG���q����7W�Z��|�)� r�s�t�A�N#ji�<Rbv�r@����ଌX��.I䌔�5�^+��/G��F�w1���,�<O��Knp�@G�4�B_�[�k�·j�H[����#W�n䐢R>D��H?F��&j�pFc[�5ˑ�/��:j<ҥ5_v)�C�kLRXT�K踰H\��~�M",���'��D�/�����u�������cN^�2���[&�Ҥ��&�tFwq��ah�Vq�.zY�e��٬�Z�M`g+�ܴ�r"�\�Hc��y+2um�������Jبjl7��:y�q�5�v�r�U��i	o����U��K4�pg�#�{s�fp���d�u������$��8	*	�8�G�t���s��=NG1ǉ[l3���$\�y �Q_�4��ƅL�&���(1��]�H�B������PD���kF�.L:U�.+����;%ATB���5%�p�3�`٬R�[�>������:�f��&
�{����� 7�AC���}�G�o�Z�#��It(�{mv��(��F��s��{{�W�4�z;�c�U;�B��z���vzWkd�{����F�᝝���}*�n�pe�Ӌ n�;�-�f0�v��y|��?+1<SI�}!	��	y�=s�r;	N�-F.a��loן��"E	�X�#���Y�{��H��B���+��(p[���P��ɚ�/�>�
�u7\���/��v�ٖ&�qc�����4���Q�I7��\���+�@b�ϟ"���&�����s�JbԼ�X�ҟ���{���u�)��p�7�.H�:[�u�BωIAZ̥
�y��HtJ��`�;�L�,�zC���?L�;�|>[��b�H��N?'��LOk�\X�T�ߐ��.b�ÅQ��F���e�s���X5C �̼D�Ã��4
Ð�)�
c�3�`#=�,�ߋc��=���0�q��\�v�9sd��"�V�iLw�Hj��ݹ� �:���3��6�y�z�RC�M.$Y����T���c"K������vo�j�0Z��b��Fs��8[����M�GUl�;��34��ˉ����㰸mh��э<8��k���(�iBgW�C	��
B�ĩV��J�p�%y_(�/���jՏ�)�����W2�����u�p[��G���8(ȹL��:+7o��0N��~b��u�-�=hs��jU���5�;�����e�L� pC�ŵ�����2��g�3���U4��&%#��-�δ��*<9ȶh��
�������SČ�#��m�Y�9�������PTy�ghR
J��㘸�an
IsѦ��Q�].r������{�E��k��)�8���\���D>����P�b2��k�{}ޙ#�j�vWB�,����J#��Z<;����8�Pv+����q+�6��_�	��B���S�;S�`��i	"|WC[�[Hi+lƥ�vϤ�K��>�I�2�4Y�zD7���z+������#���p�Yn���������E�uN�ɮ����
�m��
����bI����Gk�<�x���[*�jl?�ZO�.�⏛Q�a�0'c]h��� ��U��M�`�.�t@
d}���=�B�r���i(q!v̦nt#���U
/E�=g7V�g�_CkB�6q�hU:�z����3���"ƚj��zr�M�=��xĈ���𑗀�G9sɼp*�oT3�!e]��c5�"
��AW�8U�#|���ċ�__��,�������m+���|��:��a����c_��nl��E
\!+��~!�b(x
�'�Re�]x+t���l?;%������2�G��`�"���s1���˹��i�ˆk���17w�?O �器w�ν4�^���ŏ�o����:A�>�Ov^Q��=�ǒ���{�d����o-�p|�\^���"�n�H5��Z�kki�gb�IdT�I�+[ ������Xp���O"�?n���ɰYT �8�}�"Xխ�h=pA�&��m�| �?�(���� ��B��ѯC'�����H,О?˵ �yw�X"���wYj:�҇0��K���e�����	�#���w�TrWQ2O��:�0��³�>�F�e߄���꣌c'����u���(?�#�=������/���Z�:;�������k�%���R�s����A��!�8q�o8���t�T��L��roh	�h?��y�V�߹�2$i�x��=��A�Nn2�	�@��`�
�ݍ��!���Drt���xWd����?�Z�1��X��uh�+[P0�X���5��,^tdZ��
 a�C���R:�_���5�4���r��-'�.?}�qC,���9��c~�25�6-�X�D�OhE{0F�C��~B�q�f���4�G9?�Ar��"�s�<�9ϯi�����22�'7��`�a��7+�g Z�(�E'���-�DA#��6X-�}�� �!F;R��9#�22�ե��D�[�5�w��;����;1������2f�a��DPU�%Ho-�1�ˠB�56][9Q����h�
�gq 7V�gD㚴?�5���>�Ķ�#��`n�BpEE�����%�Z�P�A��h�lx��9����G6�󮧪wP�>U���n>0����:n.1H	5�?�?����o �ɳ���Ҿ����z��k�%ʌ�qWI�*sz1/)7�cC�AߧZƺF��d�!���8Ӣ���?�:�y��賀U5���*�v
���ڻ�/u��������*� �#p�)�4�XbY፛%򶠢*�,F�~.�+5����JB}�qʣD��<>�b�VWmϴ�ZŘ"��b����P՛��̷�l!�R�u|AX���q�4 O�O� (-�q�Q�}���C���db�R(�O�Xx�#i:`$��Y��Ov���XM͍V {�+	ŔZ�b��YK�U+}�������wF@���������Ќ��(�p��H}��L���:K??˺54?�ݷW��)"�����U�b��qr�����E�6�$���o�@�ו%�� /���t��f����q��OG)�ڰSF���-܃p��e�ի���{g��#?7��6Z��F<A��`%�������db���}�5vB�;ek|����}�Yr�c	��(��R��C�/������'{�����-]Ja_9F�	���G,$�¸#iaQK����L��ZCH8^�h�-��qz<�{mv6u�l�s��7�ܷ�7�$��ϧ�Q�zOn��2�*�j�sJ�X��|�����ޥ�������lEq��$���A�j�;�'�96���>�������zJ=�����5�g�Y�Y&xK�g5=�"��N��;����-��A�	�TN�y!���HÂ-Os��A�Mzj��;���~��&(�QE�0;I��n�^�;���9�Z~>o��^�U��~��Ƴ��n��������<.��Ų��&��� �B�Z>+�9�B�������F�����ڂq�̆�H�"�����p|��.q�(��g9�$*ۨγ����<�x��]@��ܼ��7���x-j�b׃�N�יυ�����Ru�`g�P&;��{s�CRF*��HY���, 7$�P�&�!�t�C�t�үǳ���/��`N���m=�m��OҺ�2wS��w��_ҮA�C��)�c�?|�œ�9��nO���I�D�@�2�w�v.�yϠ�GV����g*8h���8����}����U�����U��ޏ����P�r�{� �GM�1�ﯛ�e��W�xR[���ݐj�MPT柍�	�7{Ů4}��i�Cµ���Ϯ} ��e;��� i��$�g§-WPfg&Ǭ׆dc�D<c�3���;#��r�u�	�ƽ߉��֘��G��@8OA�C],zI�%�(c�x:�Uqc��*Ε,T�[����l�<�<t��;�Yt�ʯ�I�̓�a;�"x�V�M'��ER|-E7�:��bѻMW���+�?�f�͞D��<C^-�ͽ�A��Y��E(!�� S�wʪ�*�pz�R�G��.�]n��,*�V�불_[�ｩ�;*�ԊDD��9�j~�GB`�h�ՠ^w��S�`
�,� �4��ӳ��P��4(�X	~�W�6Y�\�߫�G�h�J$!��Rv��H2gp�b����LR���/�Q�NE޺��3�Y;>�ibay|p�S5�M8E�E�}�r6x�U*1�R�$��5[y�0x@/o *���T��t�B����o�%gkʞ��l��;!-�\k��ko��Aj!m�
ͦ}��0�����S�q���e���>o�8�%���9���w}�Dv�3��)h� �#8�J8j̡�q��?�h��K*��\�S-�R�D<̐~��g����!�X�/X|'z������	�����)�5 BvN
]Hb���(���%�r� �W�֟���I��� o��e
�v�^�[�㚵\��?'�^/%�_8��ˊ7RS���D��� C�Q$Y�\<�^�*`tO��e�'0Q�������E���N_����+ψ���8�#��]]���6=]_��I�LL�V1Ъ�â���:������֖��&ȷ�^��v��p�M�bO�|����«9ؔJ��z�[6�$����L9��[�L&�^?��E|��{��1�c��A5�����S����N�ؔ>�D�_�Y	?26�Z��f���92�ig���+�= m��o#F�|�;	>��<�+��c����wo��Ԧ�<B?�\M@��ygh(�l����Y�$fj�z<7�e�e�3��S�C�w�D3�m���a(G�n ��*�q�d���X�4rl�.Y,"����,[�_Z���֛�׫#��?�ig1i��|���aH�����l��n�Os�01������m����F~��Hq�8��fe�|8E�.H�8�5�+���Ӿ>���:~XzKԆ,��n�	�؆y!�walj����ٰ}3HQY^N��_(5�.�R�8D���_X��B��u�����Be����n���D;��S��6��mCUB?S�W?�z�L,3�ޜn�q&�2����@��a^�>�����YDU2*�T5�uF�����{���g9�TI4�.1�5���=��S�i5�fG�	
g�'8�6�C?��6��im�'�0��^�Fy\`�Xu52�*�"}y&#�/��*�T{�\N66TR���\8�f��dj���yg�ˌ	�DƆ}�P�IM!$aASF�Z
��v�`/:�EI��Ru��5߸]�������f��Q����g&fov��>��瀲a"��J��U.�HY�������Pg�曻m�%�l|v�������|�y��j��LF�~q��I����+gL��|WC�6i���u�����h������Bk���M8��cRl[�/
i���(�,��*��]�5���D�˿o0�o�ڌ4,
s�z��}hp`Ư��y����<,��y�tP���_�b@���;��ܝ���]b�ׅ�����Y	�2�L����w��8�i��Uw ��5���o?AɷI9?߆��A}�ݾ��6��	�W�� `5Yc;z\i;���P\�S[��	��H4-�������4
T��\M����4 ����E���R��fM �WM�wE�{�jl�C���+����q�`^Eu�BJ�$��%o��rP	<Y#����t◘�����lc$������vV�:J�)mF�5���"���FkWM�܋"Lꩾ_@�}{���z��r�;C�Jd#O�$�۔�S��'X��t
)'A(L叶�4�ˡ?f���I[ñ�����47�%3Ƃ�)��%����J�"7���v[Yj<b�����K�7+�����T�a	�
4�V�H�4��p���'cJ)b��|G�>�?g�ԂS�l�9y��s�,|gH2%�Yv�K\CtW��c�R0����MUŢ�6�q�C�WI�;�*�Bh�7U��;b�2_��Q~�
4�n�� n.��D���m��`;�Fop��&��/Oy��� �tS��eF���7����{o�՞�Lgzϸt����}s#G�w���j�߾j#����Ȣ\��ػ[D{�-�
Ԇ��7Z�fd�smo�=i�=���҅���~�U���uO� �*��`4�,�%<����c�pХ���<�E������, ��Dp,�m��ۯIܪ�~��[���X{�x����	��pb���;�UP/���W�6�Q6	��z��g-��?3��$@���A0@��_�d̹�h��"�L����ʐ�qi���mBzCrH�x:_0E��}3 �nݜ���?�w����=�^,i���F�sAЌ�j�i"a)5�� y9�����+��p掉��7*M&��q��6s.�r�)NԼ�S�!�XԀ���� ������lg��uX p(��s�x�	����-�^��%-���m]�R�%<�$ҹ��� ����\�&?�Pϲ���Τ�tt|G��	};h�P��n^:���Yi�F�@?)mD6V�(�߸�F\�U�������B+�Y$�[�W�J���K�5�jG�k'�xf�e��w�7LJna��A�S��0�G0�(����i�p��w0�:~#Ac���DjG�e9Ed�W(� ��FpG�`�[��ٚ��"�$��;�z}��Gwd��[px����ƙ��R<ڈ2���E�P��|qժ���*�gb���u�m����7����̟#�B4/�ȩDs*!Λ��������K��X�ESۿb,�Rw�)(���ڴ�`Jʼq��Q&AF�'�
ŧ��%��t��b&�f���� �C8��B(C�QE��&�.L�
�����De�;��������p�C��6�˽��)&㯀��؟�gHk���>��e���̃|�BX�f�m�P�A}��% g��o�zن>� ��;߃߄*�m5�1��#�h����E7Oէ!�O�������-�u��f��M��DI�JY��\n�Z:׈g�
�1���SK)䳇�*��[ݛ7�&�����!3�����=��������d�����_����M/��WI��N����w@w���y��V��CJ��~�����ݯ�+�<.��q2�y�!"GvG}z�7��Hs�%����y�֩r8��ȇ�?���	*6�
Ƹ}��d���9ҧ�'۸_2�L�\w(����B�xG�$��̨L|�u�m*ۍ?;���2Ӷգ,�݀R��L��d[3���$z]��	a7Y_��5ؾ���c�I6�`��"DZz������b����[��Lr��P�4��I�iy��T���\��p]@$Ame����%��Aj�D;�F4W�|n�(0\1�Z$��{5ַF���h�����S�k�:ٲ��P��ܧ�c�# *�X
�j8��!�Z�Ec�����p��,%��R!o�M�f�X�~#��~�}��/W�����"�t��b�����@&�����9��c^de5�"h@�����^e��ր^N\
��g��T��Pސ>��!�?��S�ʽ��j��q�$/��7���K� @�Z�~�$�'=�Û=��b�1T�f)՞mB�$���ؤ�4�f�Қ�!Um��C��Kn>�j��A�1|aK����mh�����;�k#��>�L0�1�� ��i�y�{�%�%�k�N]�}���$B����+lZy�`ܳ��Z"aJ�_�t��rCY7�-�-�_�@�O"յ*NYJc��۸�ӭs^縋���g��[���?�E�)�:�C��$7IIx��,���b8���c 	'��0�3��'�ˇ=�(��s�̮�ˇ�L�*�������<�Ͼ�����˓�����I#ӑr(\�^�;!�|ӷc����&��rK$�]u6;���YcXq�w;ov':�~��u�I^z/��R�q�*-�ՌM���L���÷��,r������.�ʭ��lƝ�}�I�S�`�������
��Pk�1 ��]�3�fb
�(j�����l�jFXʡ-D{?�_�g'	�;>�6G�k��!Wr7F�,v�Cu��g~/o��O���
��n�\���t�*��#�v�`X�5&<Q�D�}��A��AO�{h9�:��FZI9{�Ar���<���@C���pn��[�|	fٱ�g��-Rłi�T�����g,��6j��to�V.pe����v#S2~Guo�D����kQ2���F�)�㒾���I���j���|�lH�.b�cBF��N%S�
��d��ɯ�?��:ܲ���p:_j暀��V ��,4L�먣����j��'��[���,g[��'n�w�L�h`�̅�C:T%l;wj�4�}��M��0��o�������l#�ϖ���M+DUȂs�k�1��A2i7.❈H��b����HYFÕ��H��;�*�$�|�a����8G{�'N�QA5�� P�V!+�S�H�;-�)b�^k�^�Zߝ����IL�ؙGJ����u���r�\�u�-������e���FAsFzk%(����C�UI5�_��.Y�aw�������B{��ۀ*Y�f"����F�h�L%���&�"7�E!�؞�����rSdZt�7Vb�0���S8aI�Q0Qz�'�����tliW F>v!�?�1�|@jR5t�"��Xx�o�tNO稉y.��s�>����Ɇ���gPXsiH]W W)��ƭ���Q���C��\�(�wi?���Ӹ�no�+͚�eͶ���*��)��<�3m]�5W̿P��l��4,�^9��>��^|�1��x0��Vj�`����_jr�<�������{�?sc�}I8�A ����g�K�שF��msyf��a�+�tm�M��֥@�D=�k4v��Z]�Z dgvˍwգr�=��r�Rd�%�j�g��t^�r}���qː�*̗[��#t˶9��1>1ȁ2���Rg��	3��7E�zq_�L�2��/�s����cu�SY�N󐟕��Udr�,�F�K0�T�xH�C�(�ޓ� S���}lyVjT���tD	)�м����I�������xk#�̭�^������]`��H���NɶD����͗5�1J��밨��enA��&RK