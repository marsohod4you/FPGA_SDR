��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��pǾE(
'�|\4��~�A
��&'�5N~�v��N���Ig$($*���%m5_�3&f&�����9U�zEL�rj���K\�u��tbQ���dFr �Ӫp�;$1��p���+������\���x�,�0Vz��]͐.$D=MND�R�{d
�P=\�[\6P����c���u ��ƕ������cUb�/�{H��bI��p�fBr����x~h�۹����^���m�pjd�]��~x����x����1�`z�(O`�W&C�:��El�y-`{6��3K��9�h�m�c.hO��,f���KC�E�����O}�qSY�:î����w�O���F�$�� ]��^<���'1����tc�Ac����0�-}��{�	����������޴=�Xa9D��N˾JOZl��Y5,b��/:	�l�~}�9�J���v���v3��hG�DM�<�ol��W�V�6DEB�K�1�T5G��d[]����$z��ݠO�ߣ��ǡ�y \�ă����o.������EJE���E/U�F�+BP�>�O�=a������{�`�J����}�uk���(x�|�:��>K���@���g�9 ������`�1 ,����6�S&	T�Vl�ڿLЏvdK7�67tE�z��{v|%b����w�5=Q�"�mQ�9�JX�3�'F�;�lDm�Fv-\��T{C�x�咋䵂�V8/
��Ml�g�뱭N�BЏ|v�V1i�5�K���h(���	U#MҫG��c��N��.}�����^j��֗�<;u0�[��чv��DAu��HgX�N~�I��E߹S|{\K�g��n�����|s�J)�]d����ęBBoP���"z����`�bI��F��X�~PÆ~�U��B8U|�ZWU]˾n��ģX�ɟ��*���\1�EC֥W���{�~L��Z��Bs2�[��	�+��<������Q 
�Йh?��K˭<e)ܖ�����R��ז��?��6F���8�� x�q��r�)Ֆ��x�0���;�"������`˟I��{%SC�p�|' 1]*��r;�9b�x�:C�8��R���j+W�o~�Y�����h�U��ʟ��r�8O�g�읭L���5�j�v�e����o��C��8�R��Z��f���O9[�� �T����١�Eױd����֕O%iĊ+��>���2�2��"�� :G<�!�	:m~g>��z�w������$[���|�=u�W`�� +������))4(q���G'�7,�Đ�N�ϲ�ބ�֭o�@�ZDw�%/��E�a$���m2q?��W�0�[��*~���9Ҍ����]�T��0d{q�J��$"P���n�6���Q=�e���x�<�K5��f�?!�\L��x��\�G����{�O��L��v,i-�����\�&��-���g���j��?��������)����~&9�p�n;l�M�c��X:�>t v�Dl�H) l�W����9a�_Xe�kl9i�"G����wTw8�'���^Jk/�.�����������u��
�L˜���A}�xu��[��_a#J�������gV_�i��5���˷�AVy(��=��Ew�&�ǃ/U�'���<�{:D�����������k���H��3��{�ps6��<�j�KO�#�6���.�wʁ9'�?Fj�'��3G&��S�^S��g�.+=#V�~O�O����Y��ٻ+����� ��s��\�58s��m�Y���x#�d5�3\Etz6�{ΜC?�7����"�@����=�pw��Ue�r�����K<���
� $B��ƻ�
:��'lMM�*� �%��f��J�f��!��S�w�|�����(�#�݊[�����lm���� �:A^۶ať��4t����q"P!f���h붖��D�$�Ram�p����`��=?��* $�'~�1M�9��~����9a�42Ex,����c���$���^ײ�� 2Y�)����[�}%����r���[OX�Y�g�,V�N4\ogS���H7�-5��CX,���<�a�^~��lĶ�Ĕ��:t���z�����7�;�5#?$ħ�Q��<Z����Q�F�����i��e��W#X�'�'��d�'J��b�jJ��ʍ�&���-r�2�e�d>ДM�U���\��H�'^���h�	���Xd*�j��~j$��D��}��P���Ŭ�7���P�?�)����."��Q4m`�X��{z��
Uέ�	ed£�ҵww*�)i/	���,����x��#e�V����9�� ��v�ԅ@� a�W��>v����ݐ��%+7E726�έ?|#e�Ǩ��`ɠ�M&YqT�F�y��
'��JKq��\g���Y�N�0���xm�z��rdGm�Q5.�e5���d�����zޡϜn��7�f�(o7޾�)�ۛt^w�椦��x]��BPN�ҁ��m��;�Q	Z���y�b��ƥ{nJ�"��чa�u���t9 e�{� ���oqy>���`�]�HU���Īt����J;:Ht�P����q����V��V8��ka5B'����H�7}Z��
����\��oT�q�Ho��`���O�����%p�� �1S�5�ع��D�ж#� щI�N��V�_�nʐ=�k�����$��6<>��L;I�d*��p�k	�⫻$�5�ς���CRLw�[>���S�ȡ	�mDn���U~�{���U���f���/2�L��̙��Z�)��d>��KK�	��ˈ�|�+�Oq���%ׁ�2Q�q�ٶ|~����1p~z��k�qnM�?s���|6g۔7�Qs(�Q�zW�J���(>AVt�с˖�
�.���l߄�y�d��?��0�C4��OH��r/}7_�M(�������`�7g�M|Ŀ!����i߂����124�X�aR3i� L����A��*�dS*7�C-e5� �7mJ���g�0�{�24��*���~Y	U���@�	C*zwx�+�jO�aSp�����*�����r��P���,X{S:�sd&CW��6��
�&f��
p��WA�*���RXI������yM�e�{��V��3�|�h�
!�Б��I9�<���	�D0��Q��VJ�ާ��M��B