��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �����7��vc7 �pz-�0����)�|�>�Fu��a�&�sams�#���1��^�c���fFk�Ki7�#s
2zJ��9���

{�^�
\D��-�J���,v�O����e��B���?G+C�w��Z�$�+�ī#~H�f̳�H�Gtn��e8���9�ó��3u�1Ӿ5���L��j(':�G��^Yz	`�����R��Gf�@����}�P��GC,�Y��/=G�^Y^���y��~�=���L�7l$)d��c�7����L���ި��'�L �c�̈́��0��X�#i�(�:��B)<��JCVr�|�Y�rݽ��;J��_�=YW�H�����M֊h�J[��-2+�n'NL��|�T�,8���D|c���aV�� �8�x�wC>�����6���}�b#G�=m����?TP��Z�:5GH�㐜*�Kٛ`�S8����d���Ŵ�Vi+7��sC�L?ϫ
�x<�=0��h�}ЛZ�P���r���!1Jig��%&�0��R��8h�|bg3��(c���zJY��ӹ�=A����<q+%����
�?Β�nE+�g����~_Y�����ާ��=�
:'B��@�Ô2ӓ6�N֚�M[�j��A�J�i+���SNSjk��T"�[�e�E/��Q�Af�����t�a���ɞ�~6Pվ�2W��i�X��-�5k4Lt�MM��_�,K�S�R�"���Z&8�ɚ]�ƽ��*}� �g��Mև�%��u�Q�D+�r���~;vƌ�VП|	|;ȍ��g�9�,�k�/BR�3s�p�ٽ�9uP1P��~�����*ɫ�Ѣf����-LC���M����9�ٽ��W�/Ĳ��-�`%]���X�P�|e��И6�Gp��?�o���ݵ�V�+c��F8JI�54{�H�2z�����󛃃ӟOK<�C�NC{��!���L�TA��-� ��d ���E*J4R	S����?k*UV:�Q����[U֧������v�Fu
h����Z�3|0�\� ����mI�ȯ��"SJ�-�fWkw\"#�T��ቸ�T��r���3�	sWTrN0��+ϕ�6�;��"�x1��4M;R)^���0����_˒��N� ƥ��gM���i*'�tKb=SBK�Sk+��|�t^t`�Kz�P����,+9���x�M���B��:Z�x=7U�ғY0&�O�����}g4�&�ٲ�5젺��hM;��e�ἕ�}���)����ѳG���(�ͽPA���9�!��h�x�Y%V��<R[Œ��f��D/MlLX��;ܘف�g
��`�fb\V��P�u��\:a@�W�90�T�MU��Z�&u&�ک�]ݤ���}�	-+*gi��:�-��=`����q�J����'��Y̵�<�4l�®mA����ٶ�X�~n�y�ϧ��M��u+��� ��%r�ynw$�x]�	T:� *ES>f���|�B�7U[��s�O������@,j��,�/�NI��GC���'Ӡ�&�������s&W�R��{>��@b���_�/�� ��ɣ\�7L���E��S�n�w��8W���V���g$�l���έ�nd��#��b�^���sdc���;�HT��u�uW�*���W����}�=ݿ�%��{m�<{M���.��o�4���Vo�'�оyQ@o�V��O11�}$(TR����B�w�.�������b'R��𺤖|h���=$�q6��u�|�$T�i���y���̙��fa[��t��������	�E�8z���r����]��n�=���� $��Fu�����{HX��b�Ѕ�e���m
�s&ַ�Ԟ�\5�#����pW]�ᮒ7k]B��������z��
x�7�j�,ß�o��6[���y�EF�+H�R�D��z/+D<�{}Fr�m��mnȔ��coLe:<�T��S�l>������a�������&�9z�����X�ƭk<;!;����۞�2|��ٞj�����T$ʠ�D��t{VM2y�����s�)�R�*�f�N�<Ep3$�.�9�C��*���R8�i����{m%k
����O�h4k#���,�x�� ���ik���G�k�)ج��nZ������n�vJ�P!�~JU ݧήQ.���hi���\�}J$��˱�M�(TЫ����j����7�؟���˭e11�τJҳ�q�����
+�BE���D�dYA���b�4kh�t:�s]{C0.�Qu����o�2�~nb��7W$4�Q���ĉ���^m�B��e�o3����L7xR�VU�++����U�G�����)}����p4�;�أ��_��F��]�(���v|\p�d!t���b"�]��N_<AW���>n b�	�<SP���#��߽4��9�ɵ�,�L�a��OG

ChE��;s�Huf_�I,��f ��O�CK�	��?A�Q8n5���#� rU�@�"�l|�o5P�o�u�b1�2�zVg�?�c�����/�n�v�RSZl��J�+�����ak��d�Ե���?�41�I���Ҳہ�gu�-�Iq�#歄��̦���"�5�r�3�	]F�� MusB6�uŏZ�#������X*��k=�Ag���ڈC�>4�cH�kލo��L�e�W`Xx�ǹR9�f�m{QJ#�&����t`U�2&]�L7�pzs�YL����}8�����TH߹E�GS��F9%A�?��v!�I���~C�,Y� %���{ ��@��M����?3�U��c��9\�n0VA���<`�]w� �	��D�̲�Gu�}OSսZ�u@p�PO��91Zq���`XK�M�4������Jo/<?��M�b�­W�����V'T��t�`"��=�-FJ�bI�����^J��7�7!��c-�9�`9��������}!%k���NDEľ,�S�*2����(d�\�?�E	�|��8W}݇���ʸ'Zn� 6��`�W��Z�d�������D?g�ƸI[����Hz���'��C6�/݃�/AM���w����/��`��K��sS��M�K��`%���n�Ӿ�('x����Ü|s�s	^R(i��ꢛ�g�����w�il�b���D�\��N,.�F����(��%��^��U��ő_�dD*m,����<x��������P�����4I$���ϴ��r���$LHe�x�����}�cǿ0�KL�W��F�'����
��pw�\;�܅=�����y�
m'��{d��g0�ǻ�����"��[1��%�'%b�\�"a�"��m�"�|)�bzL.Sk]k�	�N��������k��y.�Q��C��u�. �--tJp_+hD��c��lVʹ�Jt�t�����P]�ݟ-+� ���*�2�i��" �y�b��wS+5`r��y�]��!U�G����} ��{�P�"S�ٛ!��<?)�')����Q�-�W$g�ZR�^T�	S�KB��NT+�F��I�-TA1����ڶfW>n�ٲ2`��L5{�Ɠ�*r�I��e��@pȦGe�s��]�`)/�����oC)t�CfI���[�I�"���O#X��;R �W�w����jm�4�$@���Nk�6��L}o �����ѹ?�����X<�\��|����Q/��)s�' Ħ^������Z��`��K��`yP���?��%��P�2��+�$��	�J�:`�/����e����R��p駠A�c)/�rG��Ay��pʑw��p1?�u[�2��Ҿ*KMD�?u���MVF���d���RHNJ��H1��x�G��⬠��#<{9�\����
����΃EZ΢B2⌺v��d�Ć���g1�����e���M\ݦ�1{J�0�?51�'�۟H2U���l������D�2�e����
J���\����L���>]��ƍ�V����2h=6�[8���5x��-?�I���!����L�d=c��I㽩�G�.��V���ᣌ@�<bb̞�q�������m�S�ӳJܮ�d�1��V
P�}Z)��|��!�
��E���Ŝ�^��{�ۭ`
NQc�K+̆�
��J�]�W��3
c[ǡadV�a�Wtl��}�$Q�'�����魳�|(����z�������.���j�K0���WY��E���zȱ�*s�]uc�s>��~�w��h���)S����kh��9֣u��{d�sHK����ҵ�N[���4t�mċ�n�E��+NG�����/�\�~K[r"t�G��o��U��/��T�Yf�[
	�ro�G�A��]��}-n1�榄�9C\��N��ә�0�������٪�	�ϟ.�)�#����㧎�N4�bڻ��������`a����Ȥ%H�������O���| �u���$f0�$��1{C&mVT`���8q�[4c��V�2S;�&���%��]������᠔��VՌ��t����|"�CIT{k�?Rk���R�7-�\�C�]J���R�]�Z�i`b�%�_�E!�lǗɶ_E��Oφ�,�RE]��u�m�;v"\c;��t��q;��Ac��W�����pX^I��.pl4k�{�/�U_�
:�:�ߖ@�����~�=��/%�{a}p2-�����p�Ǫ�T�zei���Q)�N��>� <�r��A����(
b��w�����Q�g��R�X�D��4Ώ�?����+���hC���=��v�gr��hW$��
�b�]�������7�ݶ�\��4\�Yh,j�W�?^��.��־H
ģ��Et��o8�' Mt������o""��Jȑ�9�N��g�h�$��k� i6B��w.c*ܷ)q�k��?Eu��j�ƪ}ҭ	��9.�%�=� [�{��3<7��}0�B����1iW�!��C�����긃�u�L�o�9!���@.�y���r.$BvJ9��J�&p?�>�b���=���D�(�c�66��3�e��Y�b������k)۷`+Xr}x����胹���������>|�iy d���0G��$}������9e8W~
|:�T����K�d��
�qt9�����BO���y�uGwD�U�J�)����i�P��Z�U��3��q��RP�߿�����Jr����k�N�N�7��I��q���[{�,���>��r����L7|�d|�QX�t�iR�u591�l�������+(�NN��K"�?Uhʘk��(����Z�,�Y�����X{wY�����;�x�E�q���iЁ�=����,E�dŒ�Kpt����C�l�}~l�m5�[�R)�d�W}y�d0���'�?6�Y@ء%(���[`���~w���D���J���������Š����wv]�����<i�t.�?�v�=��1�x����5U���;f#&�ϙ�n-=(&(�e��$Q�9�E?�`�^�p��Mg��8�7� �b��p�_���Lg�d�C��d=�����Kإk7Q�ǋKw5��D��\��>gœ�_B`���{�¢T����~�%���h��{�ex�ԯX���JAvor$^G�"��Z(��|������[Mb��X�L�nC5���H�`Ն�pH�(͛I��Ƹ�
!Shʝ�����J���Rc2�F&nq���N��Hq|���=�ޑ�
{_h3�bd�߰ǃ<��	O,�!������!Qճ�H�����(V`�\*����Z�p��7��v�>rVХm;��(�敻�z����<��o�@�ǒ�ds���`�����2��[�Ô�[3�,��D�v�������jX��̋du�bd0�X��\<�]	�OU�uS	�����Nql������V�/GVxQ�i;� �D�&��xPN�n_~��}���� �$���P�q�����-���,i"���=׿�`�8����j��B���[���ڥՂ��~��,�p�mY�V��^^��'|JAP�Z����Fj|�i�D�}����lpo5����ф��Qб��)�W#1Y�IgR�r��J�&禢K���ȩ����#諺ɳ@�N��!�ft�GMx%ɷ�ePQQ[�%����39��_��;���i������Ӧ��;�*ն\�U4+-`P��_�0#�ԭ��G`�	L$8���n�"�d��s�����nB�mi:���=�S5�Ҧq/�ۼ�z�D�)�%��g\�=S���Z����X5�T.#Ҳ�u0����_���$��n�[�8��Dv�_4�D*"d!\���
H"���mq���M>�������/����Q��
l����Wcz���o��Z�y��dd�Q�d-A�-<�y[��c�]=��4h�9��Gy�D�D]��rX(��C-��Y��k�2 ������T����Yp�xrMK&ڵ �ih'.�LĦ~����'Y�������P4p<{;5���5uݟ&��ڢ�zM�wr8�*�a������h�� g8 I564�"�K��jkE
��(��SOx�}M��'��s����ؒ��|՝Ϸ5���R��R�^��m�7�c7x����Q�ü�Q�"B��"����k/f�6�6]1��(-��ф���΋
�?����4q�k��G��[#'t���:���J5I|ͻ	��V�<�H\���4�/k|ԩ�nn��E8�z��sD� �����z% ����8�i)���,r�=l9�>l��ML�J��
c�2��9_c8k�픢��Ah�F������!"'��Wp
$5g7:�$�L*L��y��?�4�߶,�^<]�2��P�8c����C��w)�ws���i�12��ڇ��%�z$������wr�hK�#S	�no!z,�r��H�h��x=.0J7~���jH1���\m�ĚGH=�Lf�P�鍳:O�2
�O,��{��z�.d�ݠx����:��Cش�e���J�J,����Du���t�iT�LJ*�G����h��Ū� xU��I�?�@z?���f#�U���+���!�y؈K:}���������̫h���=�	�.�Y�I�﭅�Y �����`�6�0��b!fc<2�	��8��l�!�����邵��E�(J�h9�mw��*�mT�����?����T�`�7���H�#d\cG�R�9�]���<5�g�m���o�N �̾�o���<ɠ<u\ �w�%�㌍߰�\�TBy{��|�u�-�(>N�2�oT$���Z�ʨP��B���c��5�<y��(a�a��'�$��^����d��o�h=Z{��4�h�A����#<��E�Gu��s����;rJ-�>!��g�P������4��g�5�M��F:NyB��_�tAi:�^�tW�B�S��eox�jj���Β��vL���ӹ���s�%���:�o��x����^'T�y�q��CYr��=�񐚄ꂪ�0@&t�9����o�̉���Qjʇ�@dY[���!
��.��96�oZF�rX�m�qϦ�p��T��P��\r��H�Jw�7/����{8�4$Ԙ�-�F��`J|�圏X[4��<�:h^w��e��$Q�=��6o�%��nIY��$�zW��Mg����n���)��_e �f��"G�s��o:����'fH�"-���(���\c6���!,�1?��1VX�I�^�R��a���Vx�o�{�*�$)�f�=�Kt4���cn̈́�E����^{���j:4�ͫo�� �:g�C-�P��w.Y�Ș�2�j�(JJ!*K �e�����&�L���~� ��2��x�T6h%t�8N�~���D�Okz�r�4*�*��䷅Kd�2�	T�8TZB���p�a�?�o�'��Ӳ�D������,xtS�<%��'�W(�x�)
�V X-J|�i���B�9l��S�=������dV�3����H>�.JEC�Oq�a+cCɥ�UI�s��!���RU����)	-PXF�=%�X�eK�c����Κ�P�\M�������VP�U��y)��5���v�5�A�>�%�󘭙�����/(,�&�n��ꚨ_	����h��=F���
�bB���U��Њ�jC!��e'�Y��N�0ϑ����邙>��WGv�ݙ=)y��fT�Tc2�vh�����))Rзc��[�鯇v2���Å$������.�≜Y�O�bt�P�jL�'��e(	`؂�����0�vl��[@,(�����������T���	�2+�&u����]R1�hP���勖o��n�\3--*O�f�
�~������:i}\�}�̒�A&��i6yT�%}��̢���4|�1����˧�x��5<�������^������=��Sm(��h$�O����������;�h&b��M��|�q�1DG�E��שv�W;P������md�}�2�e�fjx.��>~f˒�k>�kJ�w���-b��s�?������9����ɹ�0eAe���gMހ���&�5���]Y�nCû%��Q�TpٷW$�(юѺ�-N�O���(8Z���/w�A��z"٢�Zm-������Ko� [}�2m��i�}<
������s���f�����;:X	 &�V��fs7��J9"��-v�b+��0QM�p�������R�Y�M�灲���O[w?��-M�k����ȶ��"�Gʟ[aj�~�nN<��2�e8 ]S�!��gu��c��wN2�!������8��Ta�uV�oվ��6�����
�)�����HX[B*�߆�� �Fc���yY�ҧ������"�Զ~�0�i0F�F�����N����_���ug(�tу.s���R�(�b/�ϰ��je[�`�n���3�w�Q*�
�M��	#���̘L�mHXdh��U�� uP�zIf�@oJe�w��
r�rs�6W�Yd��ƅ�r{�2|��l���YU��!��g�)rB��5e�d����a�(B>;���	g�/n���dg�m��)}�[j�������ƫ��*跀���`��ڀSa�@����)S�UJb_-,=�3`M��at����P_	������3R�5��|�6-�z�������
��3`�$A��M?��U�L���묃��L��v�;>��@LY�t�����*�K�@��6�m�p�G���`]�g�Gz����g@���m#�fu*��H�~e��ꑆu���ȼ)!������k+8.C�]�{�=���z# <�YM���=�����Zð��=��'yS؊߯S3���r���R��Jr�g�ξS�d1ژjQa�-s�0ٖ�[��Eu�)#�s����#��|4b�C�Z���9���lAf�2����b|�^��p�NC�~�u��B
�Z��]2��I4cOrME�.�w[ސ��;�h��Zl�&&����-G���iץ�##�ܡ)����!���(Џ�ae�֕p&�A����l�l��f���je�Et�GW�V�:"!��E��/�����ҶQ#D�z|�pq��}�On@2���D������K�h�V��(*����������;�{m�7�#��$z/��mVR�����W2E����l�Ba�0Ev6=\�q6�Ǘ���{r����!�Q��P5����[}{+rJ}��n��yћ����aA��`'@�"_�m��+�p�v��/K��9-!�I*lti�ࢁ`ʋ�/UI�6g�pQw�"q�ig���jB9�V�U;�;m�gX��|��Gv�G��S1�Y��VV������pl�M�HW5�eڦw���$Օ�ya��OhqE��Y�Mv���Y�J&�yё�M͠�hea�tZd���8���Ζ��Z��i/v8���	=��hWVH2 ��a9��.pcb��r�����������xnn�4wG6#��=-?�Cx����Qݟ�R�ީ �*�d�@w��ԥj�#�o���]o��+��~|����\)@���eX�\��̈́��y�~5�H���<���蠞h�C�U�Q��'h,���ǢO�����3y֨�P�w{����6^cH�j�L[ů���P�M^���,��F�f
��S�75��R�h����KŻ�.l��o�>��'�N���Y�7�$r������y�wh����F�FB�8�	�w�ŉc짅�#2'*3u`��u����k��J��%�����%��Y�e�X�
_䚃�@��7Rqti!Nީ�S�څ蘐�Y����g �r=5���N,кf����N�]{+��Bv�ᷭ���c"��J{� k��D��T��؍#�o�L�3��(�N\s�;��ƕUn��#�˅sjS�>%/�s<�6�6���ͺ��q��!l�k~*>�u�io{�Y�^ 2���9������4��uhأ�E�yz5P�=�xf [ODiۻc��3�/r�K�g�Le��~_��ԥ��K�I���P¥"�z*,G���S�G~|�4~C��AuVE����^���Qw.�x��U�	v�,޼��1S�&��'�J�5�E['K�{f>UBL!��#i_��ŕ]��Ҳ�A��[�j� +P��M��U����������}�Nc�� C��T�+�ԣ1��^ɜ�r���p�W�c+�L�4�e.`p��3��y��y38�;X�E���b4�X��_*��eCx�gu��J֚n�K�C�f)Z`��eM��.Ұ(�~WB`Y�8�3���]f��)E��6(%J���ʤk�'2PK��.�N!�����wmW�͈oTd�y��G�5���nD���Yϭ��`�l޿�|��0��s��:�Er3"Q#��YdSms�	�A=�ڶ�=�7�R�Z���ن-�{�����cӦ@������A�&��z����!���B}�p��TV���T��Yq����{�S����'�r%�-�0�����P�=�c�����]�r�(����[�[���~��ų�����IJ�'�
�6��-�'����b��'���<�hy�����6��=��t��ǬG�%�c�D'."Ȁ_�K����i|�w��wZ�3nM�[;@@��6]��I��?�)9f����P��`��X:a���w���e��G�^��rx1J��<� �N86�V�j����'�f��C�����c���=6�~(�)�۔G~u�ڒ��T<wc⚱C�^����6���Ծ���t����Wz����q��$mn2�2㕄�;�W�/B^D�R���Q�U�`�������za&�g��}���D��Ó�{4�l�{����d�֔�����2Ѡk^m�8��nX[L��--}��3r�(H���R��$m��� "�oK���9�K���}U���b���L�'��6#ǃ'}	|I�?�T1����U[,���u���(,�|��(,��،?XO�X���4��a�y�tH0��R�ͅ�e�|��\�Kdt^VU���Sx����{�e�R_.MJO�3ˑ.�#K���������Xt3��Co�[?��i'F�^�v��!�u{d���&����	���y󭍚�+�C�����
b�5xAxf<�U���1\xv2��X j�,�����,,O�=0^g��B)���zK.S=] @Y����0�|Q#V�XQ������ǫlo���;o��ڶ-���0��m"9�/��s��sZ:�>���i�����4��&�AHO�������{�5`���)����õ�慨�b�e�Ш�~	�Vg�9\`��M&��+Ų��jb��Ǌo{�+�@�:��	}Z��$ܐ��T���so	�-��-��+0*6	��E�@���]�i"��qE����w��<���6��ٜڃ(���E��똾�9MO�v��܅n�C��4N�jB~7]�1K�N�C(�3��"H�Pv�5�&��R�",eU�È��({t��|f�"�P�|d�f�N���qy�S��a���J8|X�����坕4�m+J.(�M�nh������k�G�D4�-�T��N1"(y�n-ަ�d��i@�Y���úb���h�w�>a������]�o���S�lY���F��iՔ�#b;�2\b��m�'��l'&����OQ9n��jJ7�]Ӭ��<��{�QQ�G5J�͊�hK��2�3���C��۷P_׏A�t�ҪV1�c`s�+r��<�*��
�'T�HWY��Ѳ	�3:����7�M�}3U
����ә�
���ꆖ�� �k��b�ǔ=���u���g�j�d�M�߱���I�M�W�G~m�'�i0yM֗6r��d�w�%T��d/�����O�N���42��eL�f��^�WsJP��q�j��v���7�W�B��L�ߢ�6VD ��C���q�C8���LC��tR����A����x��B7V���AVsL<����Fr&�0T�D/�礡��s�d/x�Ϻ&<p��פ�ݗ�1���L&�*����Ĕd\���ej �aʟ���]HD����͉� ����ϊ�u) �P20�����M��;��)]a1�Q#)S��~=$������iV��Z�!�-��T;|+2�j�L�?�z���g4C��\	vd�?r��=,<�Lk���yM��%+����������ə9�5<��/�rCP����� �9v-X�@��m�Ă���0}ǚo[+�5g>ȪP��*�<�K�-\'���7�/OW�;�#[��!�(\ĕ7�i(���%ݲIN��t�̆6�=#�b=2�R��� z��P��F���\��2�*Jcj�O0�I�ðq1ƶ	�2��?p���1O�f���k�(vH����h�*�R갗������
��$1#jIZ���φc�no����e��KS.��c�}��Ft�8tF�����Z���� ��z���k�O�P������.���|�=��$^{��M{3�7�8_��q�ʐ�M�q���J`� p8��F��b���h��
9��]��Q�����X><7���|j���>OF��-f��
�@�i�Gny3&V�}=��mh��*`j=z�t�4�2ټ;����*��7
b��^�*�}����I�߂Ӻi���*�.ٞ�˃']��N6|mr��.�l�ڟ�H���}�5�U^��f)=��K��Ng�v�.N"GQs��X���\,�K�~/{�5 �PP$����d`�Lu��k�Z�)�BG�?v�c���=wE��C����=.�z��w�z�H����#C�y�G3�UϞ�`��ଫ�Wſ�<�g����y�{1{��/*oh��m;ǝ���s)Qy��P�^�5��Z��� �n-���C[a�F�Sz�yQ%�"����W�Z�/� ^ ��5�({�1�T8�����vH��Z�^S��t��|e)	@`
�wѭ~Sq�7̀�L�WFY	�+�L�I})��M�]"RKӁ�K�J�$�>x��
vPh=Ɵ�n��B�De�Q=��a}����q*ڋ��5V�.O�|'mm�ˏ����s��$`���_\sUb�dg���&��U	Z#Rk�벡��R]�/��z@���x�[�5Ey��pj�m�c������0�\�K�[��o�4Xi���V⻓ ��W$�]$�f�+P�>�]?��[I"?-F�+����w��Dj��*�6��cWb�`��Kgt�.o����D[M,#PC��N�<��%�P�j��D�H���������lI����X�I��.٤P�_��-���alCH�pyE'�^��R�۹63��X�#ԁHn*lEl��B�W�͉��c�Z�1x5G-b��2q��	��ͬ�}xS��������.�h�4��r���CT�f�������WKRquUV6˷� ���d��@̽������yȐj�`K�sm�7i�Rhu�e�E8��o\� �l#��z!���9yK/7T�Ӟ��s�Í�x�/��n��s����O�Pq��/�, 6���w��XSa�����p����[vrA�N��I?z࿹(�����kڢ�{[Q�2��hް1@������v�?I���	�1O.��w�j�۴� �nQ�쁟>�E`F0_E[�g�F�B����i�|h'x�ŴK�Ϳ�@��`{Eር�U�ۀ�*���6T�lN~�<�Y5�T����P�a���������X+sF�'�S����5{��?8���:��	`9�e�)���'R���a§���m@�1x+I
�]�d{�:�J�w@�B��(�Q3����"p��%2��Ty�$�e��x`ҮE��~����gY�O�+����^&?�v.����ӑ3��3�e�3���/��[0�*J���[%�~�C�y�J_nB�^W\NCߟ��!'�0�Ȳ[��8EW�������g�=5�v�)���P�_�����&�t��=�	`�9�y����m�[�pH���ޤ_8�X�r��MSy��Ӽ���d搶m�pV$�n?�W 5�V�t[�p�O"C)O�]j�y������R��ݣȺ3a��F�6e"e��2<�~"�F^sn���8@��=d=�oX�|�7����HT�E�}S���q�P��O}+X86�|�}��2j�"��q �B�d/�N_��0�����<�c��*9!l��*���4N�?)�҉"�:�<�*�j@:['�9w�H��U4�}>�Li�*�����e$
�E�%i�\��b�nU`��F�_S�8�t t�"�FA|Ԑ	�sX��<_���Yp#�p�{Ht��ն؎s�.٣}���\L2�!fl3�*�v�G�� (~�(�KPG������<��r�ͷ�e`�}�͚fc<���+���*t+���F�sք$����LR��PA��H�z�?$�f�N�A��[r��ر�&~j\m���SGhr'�s{��Ͻ�=�=q4��Rv63����D�o��C5��Wn��C��de��I�^�Q;�J��gd��im�f_|�����.ҹٚ���o�u�.g��c�ڨNf���Sdw�r�%pr&��p�cJh�+XXݯ���~T���Ū���2��J6�����/��H!�˹L0�d�SGS2F�t׉�R�:O$����2��Y�����C�;���&� Z�>\�d%�����j�EQH�p�wR�={����}��H=�.����irԏl�iZ+�G1r:l�|��ՠ��qۢ���@(z���շ�mT�w��s�9T6}��A�ݢ���]�l�T�G7��FY7���t�@����m) �����B��̬C����
�n�ȑ�������7��r���$�+�:�ʶ�%x�Pw@R1L�	�I�b�����Z'L�o���#���0x�*sפ��Ldo�!�zI�G�2��.���G�73���k�}���X�ʡ�,�wS��ed�Q:GƁJ�N��M��c�]��h�Ȉ�Kn��P6��x`��3�]�c$�4I�ޭ����'�X�]�Hw-Q&�K�-f��1�QW)�]�i�ݵ����!�G���+��=H���h��u�?�?��w�ҺH�P����L�tv����|5>�����i�N2�z �҅���B�垓�L��d�B��Z�iN��IkO��i�"L�����u���WJ�l���A�{�D_��c�ٱ%���C�Ӂ����G�#�n[x�_�[�x5�HX��8�n"�TcĖ��x�p������'ej�6�Q���V��f���� @>!r\�d���v�偔�6��7e^1�ۆq!���H-\��D��Vm#2�� 0;C%��}9��D(��Jd�Y�ϴ�Hg�Br-�)d�70�,�.�hrDj �9�Qį(�w�ͺ��������L������u���3��y��烧�g��p���CwF������ė�JC�[����?�L�BQ�	+�R�t���DO�"xbҋ�ݸUGW�Zp��#"�.X�K2�j�gb3�Q�˖n� �M�H�V� Lh�/��~XO�S���a�����rB�|�l��Zѩ����@b�t�	���;����Ѥ�)�݃4����2�1��\9ݽ��@�"�M�լݲAb�|�r�e)�JMḢ���&^�g%y�X��S���]$�b۳��'�Z�_�H8F3�ge�6)2��,�q��|(ǁ4�&�� �fd�Fq?�E͜h��c���=�E��Q�¤N�jf�?)�e����sfB��`�����NNHw&�/�������:9�ɂ)�е*u���^R�FUmp�{����`�a�- _ے���<�={���`��."l��w:ym�	�oݦ :��>N�
O�s��ﰼk�:��%H��F	�E�a������T��tue]���5<D�C.�ڒ��{�����(�P�7u���0�(���'��>���c��D�{,�ή*av���ystX�.�����ܨ:����R�p*~r�LNn/[jD#U�L��J������]��Je�)�*��<�6g���q��aL����
���i~��6��ʜ��k�k<�i� =�2��G�e���`et̳�Gf!"���b��d,_�ǿ.�x�
���$G^��{xāQ�h�G�fӴ�s���l�����Lkyb^�`���c���7�)U�g�Z�H�:����ʅ���퐢Tr�rG<rUT2�Q�����<�%vt�"�
���hJD:�	�[Z���uA�;�L3p����jn�?�Ѫt��t�k��U���]}M��ߠr�|v͍���̡KL}h�������&�s�07�Ody&���tZ��F�Y\7����%A�J7Õ��&�81�I���tV<o@z+�5�Y8����yPP���It<�_�8N(e�=����։L�u�tM��vطf�:ic
�Og(ZX�+�v+�|���-�ͷ�I̓�E�'�Q�]�ߐ[(���h��G�è���ll�I�W��_�$���+�C�Vv�F}�6]_~�������	�V�36�Mx���Ba{j���4�\����HpS0�_��Y�j�����G�8܆�ā�G��k�S�Dr��!���z�y�6���N�;]�S��X��b4�YC�UX���&���|�\F4픪�T�bF(�N��S%���Reߌ\�X
|ťvZTza�J�s�O0�<��1a�c�7��c��(?)����z���BƤz|�M��@�T����@˒��M�8(|�[��\	��gO*��rh��b�����e�!3�O�᪖,=9��c��r獿��z=\�6���d����`����g��QU(�'�X�Tz;��ɿn����	v5�g߻��J<9��e*�AN�T�Qbq������>���RY�ӱr�#璐�3d���N�$��ʆ�7 �3���.�]I�IݐܩFv	��l�%�E"��ۉ��y7C�ϊ�I{ëK�4���&����E����b'1?�#�Q;IӠ}���'{FwQ�k2y���`G�P!�j.m�
���� �λ�t����W�j��D�;�����@.��>�v�;��?h�<��T������+������^��A�rND@.4�89�4�sп�m;vB�@�¢~C�a��(�?��4����.��H��Pk���M�P�]?�T� � f/�ljR�U[���4����܌9���2�I*�h��
��Ռ�4O�Q�/��^��e�~l������X�ˋwQ��b�4��s��3�SH$�Nk���a�c��^���(f\�'�P�[	*���{^h��=�|��d3g��M��3R�׹��AHx&�uߡ�OsGb�P@	����:[%=�'�WZ37���������)M�<�m�]�Gt���G� ?ӕ��L�K����&s��K��}%�?��*��=����@
�!�Ht�!�FV^Y�{Å v���#A�y��A��}�q:�A�Ы�8G�7�yTH�0��5�O�S��_�Yļt���W�NW���X�:Q�́0!=+��*�j�W;+X�=��&-a�/�[�@J�k����6oFuNN�52�3x0!36�����׏��y������=�<Z�V���T�}3;Y����uS�i��H���
��.�A�N���e�zD�x��`�d�
��	v=���&�
�\�<x�mK���6xe�~���6z,ꇷ�'4"�;!��l,qx�$�����~q%R�NϯR
��8���<h��-KUFo���:�C�}�J�ׇ��.mU����Y��lFF74b�K��L*���t�1LGV�W��t��LvsD�e�O/�����.���j���yR�}��DS�̳u5�7|�U�90�8������gL���R �0is��gS^��4Q'x�u�q�@�:�7�+^�M������}/Ѫ�� ��u��/��pR�3K�B�m�xi�̧L���-��d
�����,���'V�|p.���XPu�>��GTeD�z/;Q����y���s���=�g{�*�	�2ae	/�Ҧ������p؝]X�\V�xd^J���zv�ʮ�
j٩7��U��*�����s�r�}o�io%3���5��f�Q};�I@f(J���
�`簃�Bd�O	��)�Ld&r��&��Ct2��K/�B<�;%�.�1��K4�X���bQ�c����Oy�zM
}�T�R�?r�C�?� �c�rw:�y���.'�����7�&�FL8L�}���䶸��hX���aКp
�� �<��=�J���'^���k�TlKd��՝�8�x�=��?��\r��B�����M�5i11ޠ��H�
�>��t۵�@ ��i4�
:/m��ڵ���+.�i�O�ퟶe�v����S�s��v��w�Y�*.'M����}!hX��𫚽��e�������:��ׇy�q ,���0�(GH"3�1u���w������6HmA�%C�N6���`#f�N�WS~4��z�q�-���H��~�k�hQE�.%gca�n`�ƢH���@$�9@�u`#k�o(T/(���/j~7��""�Ȍ�%T���\�^��P��J!���;	��i'k�Z:��>�i`�u�p+kȚ  �x7M�S���U�IidY�^K�����C����"���3��y��Pu����.�\w�@x�?F�	�t1÷o�CKN��w�R�e?��@�G��81ٯ���g��A��ΐ����~�*�x(���ļ�P�"���G+�O�X/�X�8{���7��h�Ӕ|��������SQ?e���8�(���p�^\A�n�_�I9�%�4�����6.� ����_g�-G�L�@�Ð��#�p�B9�7&�1�4��v�_���ğ1�l�3S �Xp��n�(��&��h�	��F\��с�=:Ϥ>%���O3�\vwm���w�<�`�X�ڑ)}�BU�L)��Le�EЄ���M��r�1]��>)?��	r�ֺ"Àd��z*8�Q]#����?���
��<�8's`[�*��,�F7��c�.�LF2����ɝ���)�5zSK���Wе�����3���Ji������*"eFbgm�\>B���;��T�>�,��Y��{j|S�6��:��ÔD��-_.6��q�#��^�#�W����o�J�?������<��rt2_وp�:��h�I�f��oK!��,G��w�j��5���3�*������z��J���8'gF5�Y����iw��}-����b�џF�1��Eݧ�ʜV����b|��r`j�~>�q0�\d��B��T_��X:�y��
��d`Jw�&t�,AP�xX�^�S����zQ���UMJ1fڈ�h�`3���ia]�ByP�aLԂ\�߾j#g!*恍*���;v&�X��\l:7���Z*28���g���u���D�#=1A^�#�~��<����V��u:Nhe7���K�A�K���c}��iZ�{+�4f� ڋ���$� �Хwf�֔ok?<P��@]�vW+aEFZ�Z��{�&����g��u�ū��?&'�81����-/�RNH�̣��:�J��'��3^�f{G܀�o�[�ϐWBVdy�z�B�#��b�lЉP������M��������QZ�0��a8R^��!���Z���y��|=5 ��e+cL��~�9'q#��[M�XDW8v�� ��~0�����덅g4Mi�]F�u�F�n�<���ѢRUC9�����SJ��7	8��~��+���w'���@a��r���:G����wa�p�?aU�K������A@R���+�*�ٓ��B?���΅�������e
�ţ����/�Q�.0&��9��YQ)5a)x�Y�{��e_��<�X!.�ϼ��ސ���,��{����l�O��kd�ka%ҳ5���`� m��Vm�Ey>��ci�zܸ�O/���}�-6�803; w����G���)�_R�X�9��4���ϻ�%՜(�݀F�s��w.$���>��mG��rA{(�sp��6���y�=����ĸ���E��oy�\L�Wacf���]������:n]0��0��c��G�x�֋2��Y��Č�?�ׅ�9�#��Tz��
��Sf��,�ct;J^�I;�#�~@���u��q��g�6L�X�A�j����M�@D��Z��N���k����M�w+�T�&�^��c�n�,��������_<O�Ps���M������xU��(�fK{	�>P'7���e"��s����ًͥˮ�7���Xx�� ���)�t���(5'e�g(��G��}�^c�RS�ș$�"G� @R�������������$���|�i��ԂԻ��Y�|��5gb�W=�0�*?s�
�W��mq�`���aGX�T�ʶ*��3F0h[�'6�S1��!-�fv��J
P!�:�u3���olr臥C��f�g�L�����E�0��FLX)���7v	G���y�p��b�����ՙ�%��d�,T:��]�ؚX��p�/q��,2yՆ�!t@]d8@D��Jl�y.)��w]���.h��ّK*i��9��� ���+�����/8:�����(��`��^h_����T���hۏ/�����Eg~�d���v�՞�A��0<����?�."Z��s1K]��\3sM+X�PG�T�©��"�,���d���1Dݖ�q;�]�\_���L68�hgÆ�D������/�Đ�N��r�<���9��|su�0q�͞Ⱦڹ��j��Z�5D�!�/������Zr �����K �}J�A9pQ�R�ٝ# �t����s��ՑF��d؅ƱT@�����Ǖ�>g�+�Fs�N���Z�ʻ��I�I~@���ן%�t�_��������.~v���K�#%!����T=}J/�|��~*UW���`<�ÿ����-�1���u�낿]����5n�r/N�ҕ�T�R���^_e�0��n�CS#a�Q5b�7?R��;,苸Ģ��NIW+�ӘI�0�$Z����h�~X��������qI���$ �ws�䛪M|�:ܭ԰��C�a\�>�=�3b�(��t���}3a�?��ʴ�۝O%�$�	{�"��U����M�g���RX*1.��=�,�W�������3�+'�
��=Sհ�Q��w�~ε8���W�Y�b*Βc�Th�/�Sd��'���~Iytw11,נ���w7I��[i�b�m������3L������0�ҔT���w>E�T�{{Ȅ��fQ�`�K��v�N��& �/�l�0խ��<�s����ﷁ#��;j1�Lڪ_�i~��:��*��}W7�?��ۋ�y���D�VZ��=]�?�E������Wc'A�%<E�h�/������}�� 8���YpL:Iv�V�C�r7��L���&�|7sXsg̚�����@�]ZfA}y2��	�i<��-C5�CjU7ߏv-�֢N�O�"�q|�
E���]�yR�1����	r��8�B�{��2_xT���UK�x5闃�rMƋ�ж�0�c��D4Q�gkl�3}���h�W6v���]7�'�v3��M-�t"��}�|��<��G�.�D�Ã�O.��sam?���I=)���gv������Lx�/w�q�̓"E}��u.���I/�蠼{>n�p78$p��
����9��G���쳬����@���s��.�gD�K�տ�X�GȦ��"�NB�b�xcMz� +{L_��F�]۽kv ����r�2�_���tF�"Ҿ�T� ��������v��Ck��Ɯ����je�QE��`�gpP�'�/��]��s\2g`�{���Rj)�VIwc���Q-{EOk��6�\g��ٕz�ʝ�y=�"Ի*���Af�ֻ���w��y0�Ʊ͟����3��0A;ӳ�)��#�$