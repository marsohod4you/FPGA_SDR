��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�Oo�X�=e��F�O����
��X����j�ۤ�POd�x�t��?�b�v�JZg���d�o� g���x��ki�g���h/цƴ��g$�Zjg�=�?�����J������9
7��%�r�N�q�w���zK��� Є�f�l��(����I����}��n�?�.�w��o#�k�c�����18~�_�w��L �J�Ae���U/
�|x`q��[ӁX�Q&Rc���e��)�W�M(濯Ie���$r��vl�����Ɵ�1�`]l5�3�Z?]�P,��V��T�D�x;�(��vf4��=�>9��Utχ�h:��I�m�NH���k��)���T��0���G�GG���V�	b&k��n��_ml�`����b"�s���Z�����2����J�[�n$�[�Y�R�w-iILe���)q(I�Gr��o`5]~��F�uF�l �"�����~��.��JzF����#�j�H��z.4��h�X�ē_"(�&�XnA�w�h���l9Ra�u����_�Pzl����=a>w�A�+'k�f�~�;�،O&�ړP��"�j��G��(�3S���A �[ĳ==Ŧ��-#k�K�e�IQ�|�݄70�{2O��Es)�@�b~3Y�v�q��Vl���:���#h�#}����ia5����xC���^q�Lk�a8]��+H`_N��et��^�C�\1F@�@��F}�5脓�ڸf1 �Z�� p�E��Jo���#����'�7��D�z!�T��q@�$~B�k\����W�m�]Xb�B��vf
b��}5�; [�(�sS߽��ɂuv�諛��"����iL�������|�tB��$ѿɾ2\)�����m�.I���#$ �:�\�Ƀ}[�����o鎱�M�K��}�#��rE������*�V���hO�~�й�n��a�Ψi?h�pt�m�V��f��Yz��@Ѝ�̈́�9�4#_b=w	:.���-�ɶ�!�q�Qb���p�+�ӏT�������9;3I"�a]":�*�xc'9g�S�t�h�?��?��IN6�G#u���,�ʣ�n)B�.:@���sZ�M��������DS�(p�zi�!*2N-���I����[h�b�
�j/f(�RBɣ"&�v��#���ob[��!Ѽ�sY̓k�o(�"�j����!��p��8�Һ�X��*�%����W̷0F�z����#;�%�*�.f�B�VA㹕,~�q�T��q�	��.��~!o@���]�H}�f�&NE�F-�*�5���4i�[�!G��:BPM�a	��K��D>@����� !�o�"��_/��w�Ӗ5�v~��� t��L=��k³rG�Zk�9�e>�V���|��7:
�V�t"�M�X�s�"�,;(�H�����C�NL��fndz��-@�.lB��-&Y�
��C��0:�3�b��5"���":gd�#���]j���/�4��"H@k������έq`< (j��ח�Oml�]���Dί�$?�NA�.m�r��L�
�+��w��M�Ih3��|�m�����W�+:+�I�� 6*�t�֜ci)S�����ʉ:��O(;�np�o�?1��6I|sdV*�V���Cl�C�2�L>*�B����%�����ǽ���������]�+^����Uw�+���Y�{6R{g���U���� "\j�������z�k�,��$�(�t�'@����a�İ�����t��ŧ�)bZ�����Mt�͏6uY�.z_���\,8��C��,���_���w��d
��R���Z�ʪwKK֧�
6t�ǯ=���s�l�ĸ��#Q�)����~�jK̄�.bIA� ��� �C��O[�,Q��uBBoɖ�x���$����a�Փ���ݿ�_Mdao��e�>�d�i�1�����Q�vT�t��3Y���A.�)�ba$P�j���C���}J���D�oT8���<�<�X�_��c܆���� 2������_��Y-8I��Z�7F� �ɩUE��+5���a"z�k����ح)'��o��`��Xv�j�?���s��D���s�i���qBmT��&��k��+8�<��ReA��n:�5�Y̪.cAl�l#��fi�"�<�J�t�Z�C3���x����z ċ� M�2#>���ET�(��\90�Ɩ���6N��� 9%�&��
����ef�Wσ\��e4J�������3�H�ssi81�X�%��#��'ӷ��?bJ+$�u�OF$����������*�g10}����{�gP �U�Q/�;<  ݡu�|�t�Vĥ��i1	�n��B3�|��h]c�ٻCϺ��C,��	�:�1���%�m�o��%P:˘g����r;�[��Y�ZN����' -Ul�؏����C�kK��:B��Gu�����~�1$|scj�y\;\��:�h��&Tq�[smq$���Eo��{��'J,]7Y�bU7sq��ω�g��7�"�q�s]����/����_w'�1HkR� )���0q��.���sl�� ��V� ~ 5:U�V	ӊ�?��-�,i�����놐�1R��G6��/-/f��0��I��3�	"[��J�[$vs;�
|�L�4��~��vK�8=x)�?F���?�;[��ѥh��f�/B*�[�w�? v�幠u�~��*d��K׎�Ϟ{@�t�{�-��mR�J߄v�87�7å�7�cb���yjS	
�ΐ�)��;@m�����L��g�x�Y�d��IAv��s������.�,'B@��Ғ������P@9�)�yt~�s���;�"�v�j�=�E��b�^��M���3s5�8��'���M_YH��B�EɆ1N�{Ta�k������?���vo<�O��4��8�X��r4����na��Vv�H�CM�G�j�''y��75t
�)TsׂB�&�$�{��������Z�w��F�ģ�*f�s�w�Ax:�D�b=��vQ�V�P�n�HewqƱ�����5�tO���V������<l5uc"	q3ny�:{��f}=K�m/B����;sNA��OAV�O�����>!����/��yA��	4���-�R4�p\���� ��˙��TMj�.�k�h"i�+h��d�����?% �����Wꆿ	��ie� �e3��U�~O��e�i�S�ԴI��Vp}��Y}@j�bc�i�t5�g�A6*c9�+9��~�>�f�<��	#n�B<�Q
,v�>%0�y7rR�F���Dz�L�M���ʪF�k*�	SV��I��
�Q��W�4��D�I}�))؍���.Rgvg�h�a,�]���A��c�w~�����ڕ�awy-�-��!�c�x���]�����h"���y�.3Bҟ��N.�
:�����4��z:w?L�l5w��Z�r��?��bkc�9{�u�v��ߨB��>��N$��+,���{������Q&�ؑ��r�&%o<D44tW��|�����6j�xZU�{�Z�#�XK.>	�p�|dT>Qݸ��;�S\�=!��@�I���(�DRK@>�?��; ��/W��\��|����r���ƩI.9�ܗ�
�y��Q�oլ�;j����g�'�f�4�U���o��oa���}�+
�<1S~��r@�s���FN��Ē�B��Wv�\�4=RX�"W��0�B��.�+��Y�@,$2� h ��]�)K����
�Vh��:]�����"d�G�Z��M�� *�Um�e��S�d�o�ɲ�2����z�����X�׈�Ώ$}Ϊ~�����Ʉ~����P�RrxA���=��=|N@W+�r��O����A�Y����!�Z�F���ң
W���{_���ܷ����FHn��T�R��Q�O�bJ�ǂ���6{��y�1�~#k-���&�),��	�ˉ�~{�ϵ�ad��F�J���q�SC�QWa�B�bd���5��Imӽ�<r�c7J/��R�I����c�k�گ$@uD_!�D�m���d5O�;a�b�3�7��ih1�=�����b�Fy��P����4�����_�J��t88���H����-<���w�+�{{k������!���{?C�^1s�.��`e���2*>��R���C�i> F��J�	!��:�?,aj��C?�qAH��a��O,��%`�h����,`D�?M��UrP�{![z@p�e}D8)b$y�N��_m���Bk�3a'�l0�n��.��K�ǝ��܆��
u���|a�)]I����[�ւ�3��Rs7W?z�J̜�`�-�O�)��Mc.����)\����X�SVh�����iĴ��`9��{g�qx(6q�����U*A����X5�g��H\���[|�� 6g����`�^o��l�(����1���%�W�,)�/��ӱ�)-�be�-��s�?ž��N��K�(L�"�9��-F6�\S�fmI�
��o�3�$�V=߱x��!3\��w������(�eh*���$��*CS����	6��	9L�sA�_��LβmW�U\xc�ckH)us3[�[fռR�����A��f� �-ͺ��_?���`Ҹ�7��6����Uùz:ā�N���x	Dn�PWP����o�Ld��x])�	kv�+��i���i1v92�g%�1 �������v�F2#ȩ�%Oh�3�Q�H̄����D���9�}�tO�n4N��3����e-p��������!as��_��
,F�|(N{�1�g��{.��WH�=�m��_�
�P��k2b�h�FK�m��"jd g[���Ȃ߱of�&�.va�;�����j[
����Y�Oι��9A��7u�j�#U� Mɦ���P��:FkW���Q���xD�!��f{���h��N�Co�����7Xc9OC�r2�����M��F�YX�w&MQZ���%�21�� A:���D�s�yw��%��}� o���K�������#�?KL*��`M$\T^$7�Ĵ��ܰ%-�xs�r�@8P%�v�."��m)�;\�֍h��y���n4��<��U�ۅ�T3�M>�7h2�(M�&��E]���S�D@g���wc����&:��Žf�i�ڹ��c��81�Sj��m�OJ�T��O"Cm�F����O�3�k�
"�;��R�s����� ��<U�_&�h�a�� 2R�����vn��I���s|��B�s(at�y�=k\�h���+~�'b�f�3"�к*�i�� ���\�<DſC&���9
Sؚ(�e�~@Tn�K(�Թw�=Շ�N�>��R謲ͨt�q|{�tWK���YY��5�,	+#�B����G>��X�ٶ����-Q�_�3���!"�o��`h��P���hBT���A���sT�fa�!�Υ�m�]+fj@���G
��тI'�#�1��kl�|���R]ǩ�BLyz.��(,)��Ӱ�͎HY��5�)��������j��0В��C}���P�$����0<�zqZ�7���ÿ�mJ!�*�!#�  �"��f"2��ԗ�[(qCwo�� �^�]w���8��<���gW Fs��}YK<e���_g�����,��(;+Aɇ��[��Qy��1V�C����� "a?�����,@��~�jߺ�|���p7#��5
�Tߙ9�"B��#Rv(7�hY�o/5tG���@�-=O�3t����x���)Ng�N��L��D������F>�����sk{��B#n ]B?Lz��B�J��1�,w�x�	o�|�+L�K,���y�4�C�,kȮ�2�AUJ�ί���BYc�n���	;�C.q�M)����E���1)���<���^fְ�B�d7�w�S 8���3F��؞A�z$H]�a�Ҡ������pB����͕�o�F㲴���MY�5 �����-L�4�����r�0)~�znVb�<sگ��rޢ̿]���H���G�cTd�R;Y�BơE��Я��h_7�F��������BSK�h��zi���J��k����1�'ÎP+� �q;΂d�"udD�����2��x!su,SS%��w?�B�+���&�b�0��t���4��ke�_G$���6ЊŲ#�e}��+����g��m]�Z��Q8�(#,�n��ԙ�����X�y��c��Կ �+4�K	�r+Ot�J&�wś���B� �w�J���߯m:�����<c��'�XEL�¬l�|�_�o^`Wf�*�g�6'N���\j�i���=d���3Ȭc�'���x�a���#����~��%�&,L�I\�Ds#s���;$'e[OS��l�H @�լ��o�@���w�����	���y먿08�\����g�	�U��J.���;�i0*�*�'������"�#�����:G�H@b"�Ac�^UP%Z�!R+����#$q�"���c:��A���J������'̉ �!�]ʰ�KK�E"f��)C����ξ�`�Tgu�JarN�{�\������_~�h�r�n.7��Z3iV1Ӕ���>��pY)�% 0�2�1�O��P���h�إ�.��ԅI�y���\�}�0q؈�Gx���ltʿ�Ԩ�Q_37�AZ/�D����� �����p�S��u{���anGHŤF~�د
�j�lqu����i�����~�}�/!����h��Q�c+��SmV�]�| �� �~v;	O�R*���sI��T�(��Dnn
!����ʅs��$z.0o����}2���3�v.Ι]9�j3T��STX�$By��k�Hʕ��քr���s�lOB�	uEnK������v��[本.'z$L��"/n���"ES�/�����\��i<i0�p�-oA�����)�m�ο^!aA��GP��{Q�+��W'�.d�<���=Y�)U�'/^��$,}�olp�f���s�ԉ��Kk�iJKbc-OT���6zfP����:2�%&2�t8�523��������6O�����n��`LJC��E�b�2:,x�@�r�E�=�FyZK���1ݏ*{�}�XNI{l����?|N���T!�,~O`K�<@v�OߴL=.Oh�䘍�.�7����Z��P��'���}���-{�T�{�U���dL��������}j�T?'��rO�CR����7