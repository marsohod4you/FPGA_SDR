��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>���q�;�;�g�?�_�q�-�m��5ʞ�œT����
��cFZ��R:�'��o�xE[�I�N���B0ˀ�2|:{4�C[�p6~��n�?�Ϳ����^:٘�!,�i�dF��<<���0������� �Z�=+C�r�.3]rܕ�u���핲���{�<bgv�x�̝(,?XN��,Z�Ag!bG�I*r�@�Y�ڐT{]k���F�B��D !%D��r_����V�}$�?�o����tS~����f+ŕ���^��R)�Dm�<�!tμ)�L_3�r����ܒ�Gپu��p+����t��q�Bg�}K��6��N�-/M�wy/'�X��4��m���� �B��To��Vtq�-v����1xƸ�����k�����4�U=��ۆ�,��
G���1��C�U싺�/�� ��9FY8�����7xH��,>�̘��&�{��"�?C��X�T�1�g�g����*�:X�_Ԯ�=kn�}x' R�g'w�T�(:���y����Jhi֛,����D������r�
�,K��jgp�@�O�)�SF�Ӵ��Ei���A�-ܲWq�[�����֒M�l%���Qw'��F8��A��:�ȷ�EИȞ�p9�@���X��"&������%���CI��X��l5�����:�>ExT�� �	��@�8l��`|&蝁�JQ��+���gf�$.Z�k��vP?1ڪ6xr��i��k/��;���D9 @��eݘ��@��)��F�0������?ӏ�����
�,ϙ�2��[R�`#�EH��OQ"I�����W�n��*���xԾ�R���@�c������UR�	�R;uY:$R�hA8\������l�u���(=��?�*nn�8��չ�;Ը��W�	�S�F";���? ����௡�,�R1��|������G0�z�F�P�h�˃�R͇o�� �J�Z��^�Пn�gNV���m�!xB�JpA��G�XUO��y�b"V�rȚ����#6�H�{rmn�z��T�B�+f�y8��=�Z�q�L0r��(��khia4�<��Z�YkJA��JP�v�1
]�]�Vj[B���p�\
�vUפ�T��g8R\ /�J�2h\D�Z������(��ŏ�`��V�a�J�},`��.l�M� g�|ewk�y$��(a�_���#@��el��(�j����P
S6"TB��Sz��k�K�~i��c��5K����o���_��M�	�Nk���D�aon�0�Xk��t��ar*�SQL�FVZ\�SuU)D�S���z�)��\CEv���Pe�{ `	���w�[���/��Z�oMI�jCp�֦��?� �~��3�Qvc�i�k���?߱�%gb�S��g�� �@�7WP�y���F	����hn-u�`P6�\I�7�c��{hH@v����v��>�^�u������6�(zݔ�_��#���1�}�p-%��P��}����J�&a��Pdp���ue�	� �K��	���D\���>]��{��`�^���=k��T��ɱDQ!2-n����t_��ط�z�zk3F���d���wDt�z[c��6��E��̫����Xcp�@��b�g�1x� L�̮ƟW��]�W[��Z6������%��#�f�3a�-Q�śU�z��F�:_��H�'=-��n/�C���l0D[�Qg�e�GBy�"(I�1!�7(y�r���O�����7�o!�*7u��$���ƄCe
��C^C�ݼ�徒���b�
���JW�v-6 4�ޏO���?��գ��M�;ۋk)8�4�#�y��NW���;p�M�`�z~Һ5��1`T�"�!�Š�B�E��?hr���(˴��h8�������3�=�eO�5��bb�8�FZ�.�*�}��8Y?a|��n�O�z��`+*orND�߰�3��\[�VnJC�NS(���A�!����bv����vw��H)'$
�{V/3F��j�
�P�(䚤v�>�rK!B��Z�v^�S�!��i���	�1�>'��ۗV{�;W��I�v�83��'<U�M�k�|_����4h?����7������{j��]����b���JҼ���b�$��,���n�y��0#{&��#�Jܤze����¾I��T3��,
^v����ᱢ�aJ-.��[n�n2��9W��;�s��E#D�H���G�;��\@� ���S�J�3^wv�P�,()�D�\Z��pV���j�����H�S��7�^ǭ}��� }w�(բn�=�RŋML�o�R��N���_c�g�������a��5{��`
K݃��wm�>�C]��%`X+�����ٳٍy��b*������|���{6��#�ҝF/g�����8~��B�1�3�y��.5�M#$��E~�4��u�fQl3��i���
���]�P��Z2iS�N�L��H�"��Y���+2�w��RB�]7��������ȏ� 3N�(�]��W��6t:�&�j��Q�,)������C+�$�>g�}E:��ѭ��0/��T[pS �x�p't��i&�1�Rz}�� rF��V�����;±:������QXe�Jy�6��������Id#�<)+WwB_%&�D�p&��[���tܹ�K���R2c�p�Ě��CQ��x������U@�W�f�����s\OǬ�Ϲe�gT RN��Eq��U'l�ѿ�O��͔�%Qga�q�ց]��9�Ǟ{���#�St猘?=d��`�T;���6�� ���)��9V��A�Q�0���{�JE�9^J]���WN�Ϲ�9u��F�+$����&��Sw���QqV
��8F��_�렠rb�eӱ�C�IY��2�}1��C�7����=؏��̾,8u��ҩ����¿h�bԿ}(�<>��9�����^�:�n�l��=,����*:|�m�L42t�d�p�F�\����$Y�89��q�"��w�9��|���j�����-�N�=?��&��c�Tg�V�Z��|lx���e�(��*��F8��X��@�?������=�K��O^���/�Ѧ���]>�U�[�{W��Sb-��c��$)���*�512դ��g�{��&�mq^�Bfܡ"�}ށ?��q8�{Q%��;�H�Ĵ�tI���J$G<,�)���aen�6�ܦ�/�9c־�:�k|!���{��Ҋ��y8a��t��#Z؛H/Ia�㗹���"?y���3���(���!0{dgbb�0�s�,��8�3Q�T��](�{�^�^�I�3��x��H�݇�Mx�hئ�<�M����5��Yq������$�U��`9����Nɳ�'U-I����ћ[zĮXJ0�޺} �	��L)8 #�x�&���P�q�u�wq�U�  :	7�������90C<Р{�����e��ô/lq���M�*��њ�~t(�*��;ֵ�O��M/}�.���1G"O;�JX�]�rO�HI��f rYq��<�{�sua�DI�����S]:����-/X
��|S�,
���C9�6N��9��/
��ER��8Ts�7ge�>����D�z���)C0÷Y������`��Q 83؆r�跂EBo��#$�[w<oM�?$�V6��g>�|�7��lF�qR�����ý��53� ��0ɶ���E��s�Wv��T�s��@��v��J�@�x�ׄ����^�4��U�]�<���pk{�c��'��c�yr�`A���9P���
�C$=�['n�ҩ]0�n�A�y6�B8}�����v��sJ��w�B�y.��W��Ԕ����j�[#)d;3��-o���Ę�����BwTs�TVR�� )!�K��?����
��L�@d�ȁ��I �Yt؟�7���?v���~�6�)'x�#�{=OT���S�&��)t���Dm�9>QT,�>���U��٣����8-���У��uP�!��l�Y_<43ۂ��?o�����/�|O|WEm�������9��_��3���u=K��k�o��v�QG��;��E�����҂�p���j��e��x�qt�o|�1A�N���|4~���m�4����!��xJ}�Bn�.��8�]P9��m�B]o-�p�i�r�Ey�_mT����}����mY��VeY��<�s�5X������~Հm��Y}���eq�S��B��oN5�KH&�ֺw����m3J�%��0�9��=��fO���zYü�ރԖ[�H7n7t��km�\s��K)nHe��HԟK�;�mo m�V0Gj�@� ��ʑXZ+�i�mN�qN2r	�� �����ˍ><}3�,�.�a�@>����p/2{��	� 3�����;�:v� c��g�pZ��$*�+���A�L�{�>�T�A�Y��-n��[��j��k��.XyS@�)�IK��{Qe���\�����?D%����}&2W$ލ7R�⟏ڳtw�Z������n�矢pmU�g�r�y|��l!�ɡ�\������)�IҘeyY��e%�_�:�@1c�Cp'<��q�O���w/���?��$8�U��S-�h����>��}�?1�;@�&q�'�	��<�e���h���`<��V*��Yw״޽��8�c���m4�H+#�X&ktM�qKa��d �����*���PG�r̫$.�v�J=O-�ȧ�K/�b��WO*�	��K-���+d�d���9]�֔|�)��+;yԴ��}b�4P�9�>q$���V�Bl��6�m�sAs��x�nX1l�6��Me���x�����"��|�d�?��u����K���}w����Ns!�^IG&y�Y�!��;���tĺ�Go+4@��;�d(���EQ>�T���H?�4����N��HD��v�z{QR��*��A\�.����s��M�g���[�?��2�Ƕ܈8�/���v³�/�����{@��#ϣ��+�̘l���1�l�F�m��US�7��0�R>�ױ�u��k�ڒy�W�͆�z��( 1�kR|�|�H~���I^�D�ئ�����C�\�x��K�}Q�Y��\B
��&eI��{��S��.� ��ƥj2�,E�&/�EF�t<�\/-�S�3��XVCG�u~�fU�����.Ȏ�?IM?(l�KS�	U��2���E_V�O��9���zO�׳߾��!J��O<�u��r����;ŉf"1[]� G�6�U�D����'ɠ��z[n�e��!��֯�/���Η�=�AvY�LDG����p��єs�>ԭ!q��5��q�}07��J��0c�Vw�"k�}=�XH���,�@��V�)�*m�<��p�l�6_P�P7�w�'I�ă�݃n0� ǁ���"��q��^F;}�����bo,��(�}% ��|]X������4���'�h�۟�禣��2���"���M=�)�(�r��л �?
�Ø)���.�����d�ӱ�
r?x��	? VS�ߵm!��}�Sw�:P"�����Tx~=7X�z��5]��6^�Gt=qY�59�;�t��E����m����*!���}�vgb�����q~�췻
?V��4���^�8����Iy�,���QH2�y';������L����7�Ӝ�Ƭ�$���)�;զI���|��%�V�;:��v}�ʸ<�i�F�~�M�H��ed��꺑$@0�u��O6G3W��qv���f�8���@_t��ņ��H[�zf/}3���V�h�ڲ'>�Al3��X9_ �e2��6�z�o;t�:n^�tYY`�} &�#.BC���_�_L@i��K�+����W�V�а��e֊O���4�{=��뎉�����c7`p0|�Y���~���2+
�]@D�P� �?��}�92K^�MW�&]n^!�D_4I´k~Y��ۢ%<��!;�mx�Q�7ǸG�1�oyQ��Ƹݮ+Ō�U$��*��l�K�-�ڊ�Y�ԍz�^�:X#�ګ�H(���R����]���gE+4/o�ܷ`���Q>�e�ݱ��"�G����������oo��ei�J�W���2�MC��1/���8���A�ɥ�X��(�y`�]}��⩲(��ͨG��sP��}�OT�M��������2Hml��&Y�?/�t[������`�T~�d��w�P�����S��[�<Ek�&�-Nڥyi� F|��)�3_%6��a5Y��7��`��ڍ��z�]<�z��8X-�$���D}"*���!H�@R��_ry�Z��(K���e�]����b�=�S� 0��'�PYm֡�����)�U�3\�f�K#��S���yb��e��
yG-�;�NV(���UC���0`�^����n4���kt���Zr����c�l?�3��F�fvT�# ǴhY�$F�][�9\̀�y�t�8�S$��e��;�}Wߞo⟅�\�զ�-'��n�j5�:��)���MS �����a�UT�8�É]��ڒcD�Ň!�&��b!ȗZ�q.^�H�m��{hvdFs��lu�v	MؤJ)�$��f�zյ5�2��:8;Sr�X^6�3�Zy��j=Fk���s�
�w�8�D�k���ܳ^Z@qlQ�/~��֐l�x�����=���Z�P�@A�_�?�| D�%�t�>(V�u��i<��X���W`q
���m����;�Ĺ�pz�$������9���`Ę��T�f4 �'�0��	1�W���l��WL>dO8��pA��M�G>��m_<5οy����`y�)Sg�f#�?E��^��
�uA�<P�Kj5mG�1Q�ᆮᮞѼ���v����u�!^�|�� f� [�8}��}կ^�ڔ)iMvO�bu�Ō��'͆�� �NB��|�OZQiCi
�����@N���j�;�խly=�����'����VE�{�>�|���#���_>L}/�W ��;k.�����#�?�w2E8��3�]3�߇�"U�=��Y~�Uc;�K����O�����Hm�6���Q��Np���
����f�r8�$��R��v�҆{4H+7J=Er��B�����H@����$>k4lB�$�u�I���h5�QBcOzǿ�
��^��4�=d�� ZG��g��͠�u(?e��iI�����Kã�Zt� �P���g�!��D=�]a,��[�bt�l�\9S�: VnQ��G��=h��r�qB������X���mb
��~GZ�ځ#qR�lw�_k�a?b-� ̭���w�}NG��$-����n�?�=c-�w�G�����zuxO�'3��8��՚~�#-])���̮x���@�;��~��V�������7`�������b�<N��'�I"
h�ԓ�al:v�%�F&뀜�Y,yľc�˂
۾{����e��w�1$m�=D��Sq��r�)�'^xS��*�]q� ӳ�2Q�5mv�tlo(��9t��ޯ]l ��L�m�����5�|��T'�m#i1�vW4hX>G{y����/c�đI��o��(�p��37��.�"?�ᮡoh"�Q"[���n+RKg�=����n�F<O���dk�0�@a�͔��ڎ��*�bq�B�m7�m�!�@��Xj+�?]oC��-���0�zr
6X�P&��P��Au��'�_�T���hY�Ƹ�x�^��'�}K�O�i_��/���u�,�կB��*f�|��F�J�)872^�eL=�Ò������ݲ�����?�s7E���~Քq�2���~@�7�9�+�������e[�Z�+��w�:�!-Q^��n�O�ػ����&$�`�Qe�MS�CAN?����1�{u�P�c�ë�A�I�rԴ���oF�k��.`�b/m1QƊ~j�S�÷k�����zu�vݑW�L޻���!�cwh|���".��a�T��ۘ�"�M�됴F�����P!�* �%��;����7Xd�oqQw�R2�R�Y���,�x+�P#PAKP<�y���)�6E���Z��B�|g�-���d� y�͔ʟ�ȋ�$.�H�)�
�0$9�(ƭ������cNWu��w�/�aH�CF��t���S�j��P�\�l�sE���{�2��Ӗ�Y�m7M���@|���}��� �"Y fA��n&�TOy,���5�J�������y�_��L�xi@ڪL�p0^ɆԈ��C�rzRE���½m*���"�Ʒ�6=
�CLs���/V�n��xⰥE�C��(��{�ܟ����	��3�h��	�ކ�V���ˋ��+j��F���D�=���S�ѱ���'\��՘���܌��w�W
`Cb=�s�p���=�����fa���%�'��6y�_G��X�r5�qLܼO���R�VX�ܥ����Ύz�`�o>ϥBS��Q�#XZ W����Sþ�М��=4���&�i��o���f
����gͧ����P��i���@��2��A�zmZ.�Uf,��I��e�D���ԃ56�t���2�n��=Ow�;;�G<���(] ���oB�_�]UpX�a��C�8����٭� p�72�5�z����W�,)�kq>�6�L�H?E�!�܆ 7���R�����J�M��A�0�	3 �۰36En��̶�t�x��\����T�ԡ�Twt��o|S�L�0Un,����[u_A^��Ԥ��$�N��z{����J��rCҽj������4��o��'1�#K�QV�%�cppx:���
�9�E!Qd��X��X�ޟ���
n'X�o#��S8�a,�R�w:��g}.��;3�9ahi���4,���=����HU�v��_,��F�I�"܍�ڸ�uf[���Ֆ���ȋ9�f5DЌ����"AOˈ$L���ɱ��/�s����I�)b�Ѫ�(=�]�C�{�D�0L��<�2��eͻց���TQb���+�I�]ڬ˓G+T�z!��J׾�H0�B/>��@nuc4io��KhZ��j!�0=��օ~��9��6W?T�lIl�v
0Ѹh�.�-�)4/�ˢQ��c�\gk�rg��x�1ĵ�7��Aa|hi�l9cuDJ��=\XHY<��Uؖ��߳b����l��tx`�;����y��z
	�If��Z�P��$h�~d�>�+�<IK�o��w���7��5��J8#��r�ۼ�ֲ"��g�K�屫tf�4@jKu]҈�%gAk��ºt�bi��J�f�u$�&n]oW7��ꦄWgO1@|1o�F�3�5�i ׆,?��P��Q�\��ֹ�9$�W�k�k�;6VH�wŽ�؆��Y�GQ�]k���rSP��Sc؈#�n��J�w#���t���9ί��3mk�4X��m�Qr;F7�T���B���~�}u�Ǔ��;���G�YR���m�!�"��
	�$�jT�3��]y���L���9�"�e��ч"� ����)�Z�@�n(=��~�PSR���R�X��W�_L��Y1JǨ�h��J��d�RF7v�[
k=e-�n��(8.��{��o����=3Kɑ��X�XB��@���(Xy�k��b�5�Z�r��C�RL���"IQ��hQK��F>�L;ƽX&1�z�&�� %�!`̷��6_�.s^ESƢ����X��
��j���y6-G\����MB
�{J���ze�S�(IX'v�~�@���5naUD^!�!�F�b`Vmeӯ>�����'�> 0G����hV�6�����jIC�Nn�4J���-Q(�[m¤�	�Yq`	��R�(�=��\�1��A��f���r��Ķ{�:��/����[w�;����+��8��h�	H�Q0iՄ�磊!�J�촏.�u��D�n�H��q�B�����xE������	��G��R5�^G^�&�e�������
贃�&>;�\�ǆ_���=��on�yͪ��i�<�i"����A��9=�u?���
A�0�\ar�ti��������=(![M:x�=/p0]��D��|�pnQm�]�@Y�&V�5^�K��
Pmj�.���TSx�ErpL&�Q٘��]�f/�WC�;��2MO]��������+�#C���b�yj�w�WSQ8j��ԓ͜�n����<�7ԐLh>��X]��Z�zc���<QO�D����,��w�Uh�*
��mÞ���h`�'�)�./HH��n�VDR��@�_N������u�A9Y.�Rs�&�͒���������Z�!I{k��Sp~z/'�U�I�NY�9[�I�u����/�§��;Y��n��"u7[҆V��8I�~S�<^�����P=a
�`[��S焠k^[���8X�q��&�e��r�S�0 �61�B�)�,�Dݣ�,Ԥ��#;�f=϶*�4�k#��	C @�/]ҡ8�#�A���z���E���7����ٰM�M��8�2�+���
ap ���:�q�#m����{�VY��
Q�s��JSܚ�#k�ڗͩ|ӕ�}M��#`�ٗ�/�$�R�?�(�%u>f����S&�.������G�o���܏޿@7���+Ov�(P,X�y�I���`���^n�m5�JD�U��4\EO�y@�"	~���*��2n"���Ծ3F֡�$�4�1�e/F�X|��F�\������:��2����M�C�Ɛ������� ���	N���s��BB��Y�^��ү.�^8
Z��&�����3�7Ccά_�Z=���d���V�e���*��ݼ��@�B�H�����N!��^ �y�� ��-Jh>�ب5�k�MG����UP�i3���Y���7$�Ret�e�g|k�V!�.��k�F���R�����JP���ĩ�ST ,y��dZ�m͈Z�Z��y�i���R�6������߉�N�Ș��^���&����MU���y>Ù
H����0��z�7�(�9;������� ��ɼ��C����VZ������:ȩ[�L��Km{J���ʎg�`�W��x5i3��.ʶ��!&n�?����ڗ��8�����Jڗ?�p�Y7�D��
��R�N/��LvV���d��͍����Hp��.e�9���P�`ݻ�y�J���>��F�g����q�����~!�s<��y*
+z~�~�3���kC�P���PĐ\�ʖc�g��rt*S��}o�y�5:��\
����3iߠ���5����|Ov������Ϙ�\���;�fpu)�z5
H]�:��Pm&�.Z�g���:_[�f��'h���F�; ��c3���b|���"��x؀�:����8l�1�Mc�7`��])�wnĳ~&1q:cz��O9j^���7�RaO3�D���W�pr��l[��H��Y0�{�r�G.-�������V�I�����ߡ3�l�kCӒ������4�E���@]ʧ�-��7�A!��̽���h�z%-������mpT���U��)��]g�gN��g}S���Ҍ�����;|�`^
?��+�R�����y5:��}�a>- N�t�?S�z�uK���{�_�J�]����c�_Cb�!��?�_�ܸ�����?_A�P׍yЅ���t����?��3�u*`}s�]<�U&�!�����^c� ����jT�|�:��;��6U���x�-� ��G!ġ�R"��WOf�A����QU��LhYSM�+�?5�Z##�6��|��M�*v��Gk�T�ګu�᚝�Xq"��`�rM�* �^�)���L��>]}�B�<�|Q�뿍�4on��!NK����`	۸�nq��"�K\ݭ?��'Xa��3}���!�E�b�8�Ca�V�U�$�ev`>8�nE��2�Wi�n���(���4@�I�e}���B���s{�{���}%��$5k�I:a�b��/!�����.+*��0�
�_����x�g��I��ʱ~�uE65D?D� �0(�|�������a�
J�-R�Ιc�� oU�)3��������ڷ!�L}i�E�N����82	Y
.;Զ�Y�l��yx��璡-R�9B�u��Ȓ�m^]�3�KA#9��^c��DX��3N�
�aj)P����hUZ%�
j+��� 1��3�f����Y(��+���[��ȇ��e�eݣFe�>o�`h�����YX�/�0%���-aٙ	��������,�?P�Ի���:��2or��g�J���O{}��C/��c�@�<��'ɿ5k��g��\Ow��Q�Ɵ]�4N�����v��s#Wv%_0�t�����,��ݣx�?�JA�,U�1�T7rF~�P�v�ڴ
dK��:r�ē�߯T�|^x����� B�892T[+����H����U�zW8g�^��{���8����L��g��a@i�,al���[Z wQ�}|u��F{$�1�"���i*�g�o`��f�q�rH��ޫ��m����]�E��=��_�J(S�-3H�7i�p27渒�g��ݪ��v��R���Đ�<� awq?���q�ᕿU���$�ɌY��L$f{�oy��N@��4���j��Ի��U)�gʷ �#[	r��<�bqS�}��m�H_���O �6'�~�r���Z)��1�gU6�ON�����������k��h�f,��R7(@�gx.\���]nI��_�V�1^o�q���'Xn�J
GS����?��rdZP��x6� J���|Q��OwP�Q������R|d#����h]�@I�;Sp��4i���D���I.��8���;�Qd�КU&�����)+qs�N@7<"MF�2-g����]�T�|����I�ہUn��}m#=��t!o����F��j