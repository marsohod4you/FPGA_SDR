��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"a5���f���wR����.F�o!��5���?���0��\�9���D�
k�A���F��ӫj�Qª1h__��m{;�%&k��i�B�h$��9f��#o;����YO7!?�:(tϷɴzw�^f#
�򕵦�ڤ$�J:e
�%�p� �=Y2g���9m�����ᨌ�)I0���m]���xP��q4�+��V���b��5�s�&o�[����Z��o�����w�d����^|'F�v����:U|�F��N�\h&.{���&��jN��� t�S���J�,�#�AI�^:��<���DY�I��uk󜊟���;Oc(y���f�B���B@7�X�__�7�N��7Qz���o�)i	=h`�R'�銇��Ɠ����w���~ɣ���tp���+N�SlJ���T���3.C��0٭�MϼO��]�2Ϧ��/�/Q�mz��|��э���B	��x�=+k&L���J��
TWJ~�Q$�`���t�e���gi���`u��Cd�_5���A.��É�!�7�*�[w,�>j�q�Y$���i��e�Z�*�pR�ٔº����_�� ����������[�s�8ȷt�J;s?0
�J�O���nj�O�����_e_J��]SF��E�0HM��,�v�!��Csd�9۸Dd޴�$�NR5Q��!��Ⱦ��!��^$eU�@9G^���7�
k�o�]G�W#�R�
t׺�Q�NM�}�0���XRـoJ(�$�s6�*�f��I���t�:t[�Kтds�\{�..���߫��7x��)�x��?��:VZeZ�La!��@��ڛlDS�^���0�D~do4i��q��?����Gjl����mM��| �3���Z�Vl��~��&��6�눻g��(5�yGV=��u�]�z�SXx�����enb+��߯7l��]r9n5�w!l��3+4�y�4z�<j�I��71E���1�
�����_���%!0�++�}V�	޽f�w�?�5LS��� ���E������ߥ��h� !ʤ������%T���f��l2 ����Qqxc �D%��K3�$��]]0���4J��.z��e*�*(���m�L�g��S�P��O�^GΚ{l����%��oT�ל����}�9u��DG�=���fi@�Zb�_�ky�u@fH�z�Ie�X���S���і�H�S�6�W&I�/�= h�ꈖ����s�_-r	$�����������ԓ3��e5�WV@r�L_
2�m�y*�]��?����/8��ޥ��Qۭ����d�{���}�����#�8�&�X->^��5�p��0.�BĖ�H��.�F�@����z�p�M�0�
��	Pkdu��!��OA��_�W!�]�n�]�H:������V��)��7�oq�,S�J�o%�W��&�0��2e�X�L|e�VW�I�g�P�����'ΒQBCʳΗ�͓xƖ����3��͍��8�ݯ������NK\`==�|�,�m՞w�'i.漶iӽ�%���^���?�{��n{�������l4`�DM���k!s�����.��?t�S|i_W�qKC�W��Z`.L�j�˸u�'�֤��A������-����
�'�H�o��E�t�7��"`B�*%��Х�&��(���a~�<���m�Hut���G�c4�}��:��_v�P5�Ⱶ��S�����Jw�C�͐.�c<B���U��pJ����4{gu��^�Oj�j���:y�TL��*C��P"`09�u_� �9�(]U��>�"�Ij�M_E���d�c{&��Z8F��+�By܂7[�aDƏ���i#v_�n���X7pb�j�:�/1�����8�"�	/L#�Ƭ%���'�w���b!GrG?6��Ǧ��A��K��M���ip����Q��C����@3V���Xg5lH�ĿL��������i���������@4�oYb�����m��	�o��G�/l�fSe�Ǜr�3�"+G�Ȥ$�-�jVv\4�7qi�`^�N��	��͂z�*t�ߜp�bI��r.x��R��P;<��2{�}��(�_�� �#yN~�"\��}��J �o_�'a�-gs� !v��q�U� d� &��~ y	�����I�%Q�\���O�t筗���C� `�屲��+�B���5.�tB6�]��x�\}J|)�7'zDL;�xP����K갸_��՛1sr������9�v-G�'��ٛE�U�2( Ң7��.�\@߽-�o���x?�W��((7%9`�6Eλ�([�I�\�+�rcb`��Y��p����J�3T�)(�?ԏ���(}X��v���G��T/J�OE�ٯ��r0�Z�$�]&���X���'O�����!\Ae#e��=����fo�h��Q���2��
"	l*���hĹ�u�ԱGi��Mqs�Y�CoL1��N���4�vƸ9���9�T�I��<�l�nÃgg�ވ���c �'��7.�n����ol2�.f�E��*��g�|�ߖl�[0/p\��oL%��g��R� �	)�zsL�J� ��47����0�~;��]v�e�@��#"CU͓lQ����*�t!r�Z�Ӊ,�E�V���>Z�# PAa/��`Y9����j)d+��n@OX���s�{�3���G$�k����n��~d�����@u��E�Aݚ��5�R�.��� ��������-��}�;��,*;ǃ.��ty���fp܅��	��EM��� VO�tk�����L!���A�_�N��u&k�R�?��(�Q�f+���0#C�_ߏ�O����8�j��)D�K��Ⓐ,��[Û�s�Y�?�O4h��[�?_T1᧒��M����<8���I�+���Ɣ&S�� ��ٌ2�E�jv��&��wvx�Pi���qjjF�A�����,�.�G�éF����{�m�8�iѮ�J���Ϗr�1��	gq4�� �Y����槵�������"?�?!��׶�g��������G�jx�����-;�}��6�;Bw4��4��Ң�L��1/|���G:���؜��>%��i�-2�FR�Pe)̭Z��VL�b��_� ��-���t�u_E�=���d�J-P����k���X��"�����M�:o�F��}!,��_=��$[?��ʰ����,-Uy������������}�b/���O	Pq[n_�uhYȓ�Rb]��|J�
QEs�-���i7w��&8�|Ԗ��"�
�Dgد<�l��QT'}�3KZ��%��e��Q�T�B��Z�"M�L�9&jA{?K� Q�ϩ�_>��5�w���r�Z@ڜHX7GA��JTp���'�d�cDr�R�SEPF5�ռ�ժp)ͣX��G�<V'�tK�<n�x��i�#�"$�5YXȓ�X����_X���!#���f/&�ʢ�� �24A���$�e�l��/
!Q�L{�H���`}�����yo[����q�ڵ������Ֆ:����� L�ߥ4V� V)0��IH�����l6ц	o��\?4L�q̬<>d[.���E�i^:�����m̏�׌r���6t�*E�F:穴�6�]p�{��Y��a�s3B�=S sej�Y�K3�:���6�@Zb���|�ݯSR������@�o��ͫ������� #d��#�S�e��&��Y�5�g�9��A�Y�Oe�bS�/�u3���	�+��9��n��p�a�eQ���ҏ,2�d���rL�MX	�z]����s}F6f;̶�Σ��e��/��q���K�f ������i%*@|�|�@�i���\��ˡƽ ��S�V_�Yr�x-�C�"��8�/�}�6K£j�%V�E���bL���I�@թ�@ivx5/��ƛYx=lQ��̠1^�ZE� ��ǚ��~XuG	�a�Ӥv?wY�Q�Z=�1�œ2���$O߄�����G�]��w��&6t�y"�^u�q��p�GW�7k�N��v��X�D�0���)g1@ni��YN���2�0�e`���M��A�hk�$�+f�8��7�a���+���K�W��8�vQ�Tǆ/�B���2�hftt���5
��L��]b�bz�����.�1|5/>V��� �����#<�l��>Y�d�s(i��,SQ]��uCٟk��#����E�pNѠ@؈=.������Hx�*��ؤp�K�;ـ��y(V�3
6����<�j�3`��c��l�L��8t�����R7�kK�ڙ�y�
����#x*/�@���sl��Y�t<*s����p��$_�a���#4Be�j�I���9��u>�����b�bK�S.$r�P��JnϜ�A�b��q�E��K=���!�P��H�����+��iO��)���)�	 =[��'�jZO=��?$5�&2�C*?j���.���̧�NI�	XD���E���u��spkj�4 ��D��K���ǥwNt6�r�6�+��r�%;����+w�`���(5|��?|��J�>Q ]��F�M������SX��t���d����`L��4mʨ�Ű�;��
-9t��Q;q��vIw��)��ԍ��_����؂���z���!���8�;�G|��sLֻ!�u��f��g�P�s^ۺ07� ��MqN�	���\7�5I#Ù��_�QX�;�����<I��C�/E4����
� @%T�w�,��0�;��}����yp�X�����;`�X/�]�O�W:y)u��ٟT�6A�|+�������������:,�������*�j��&�NJz�z{}�{��cڈq�M�M�,M�)�����������d��cͯhفY5�X�}%u��R��j�XA�E��&�H󴮸�����qs��t�`s`I?o�G(� �`'S���g��f�J��^�2E��'*�.�/��`�!P�g�� ������3I��K���\43U�{�>2Z��7GZ&`Ҽ����(ubah�y��#�X���.�0V�W��-%*V��ES��&aQIw�9ءt.`�b�#�J��:�����y5�E����cnY]Ƞ�Q~qh�F��ġ�T0��W\H���Qs2o�j2�F�hs�?����UZ�����5�p��U	�#"�,'��e���E������b�Fg$��-�t��|��2�.���ȓ%�^�Ƅ�ۼ.$�ե��a�2��{TC[8�#��
b�"x�|݅�e^&D #��Qo�f��b�7Sn�U� JR4��Q��cS7������I/��*NB9���1e�В���pb����/��/̧�Ε���g�yV��)o`�o3E�rV�s=6ab��w6ct�-�7�.�����^YY$vHh�	���!9��}m�V?����em�e��ɍ�'����hr�g,g<�ƥc�)P@���Hi�(���&k��c�s�=�lڵ&��F{r�y)c,��K����[�y���e�r�i���x:S+_�M.���g�|ʱ�x���{=��o�(_���F�������H��E�`B�N�]��w��K�4����CA��4��^$[����3Bi�ƫ�B{*����|��]mv ̱g��\,�z��vE�������2���eVt���xa���<�y����\7?�+��f�#��'�8�t.ޡ����g3�0*��ng�bh3IJ7=�[�gL��&��S��8�������Mй��޼��Y�h�+?V	��H��Li��1�e+�@$�8���+qob������(`��{�	TB-(?u��c�F���dieV�J\l�5�\O}����68|��r�n����➁�v7c�3c���K?65$�xwa�݉/x�6H7x:F"�2HpM�� w��|'�+}�h�<$"��rE�����Bq���S����J�7ߡ]p��b(.����l,�p�qWiW�æ���M`7�(�ě� c7c�K}= )![�G���%�,�	awoa�[���4�*#��+�X@;��E��p�پ�]!]̅�8�b���[qc�lTG6�ԭW��Wv$u�!�;V�%��[���Fu,̶�����"Ǽ�	YZ{��H����	Vk�� �"#�;-#֢�ق��
��<]�r܉���(�-�[�{�="ǡ�L��ɛ��a��g=zZ�I+xxS:AT6���������)�n׆��H�S|�ؾe�Ddz������n:FM�e���@��o��*�$���N.Ȕ�X�Z�<��2a'����#8�jA4��#eA&'c�sJ���E4�}��C����.J�Ur���r�y�-އ�^N����B1�T�h��P��г���3��4���Ś-b8Z@��{H���S_��>Q���~�w��?�~���2�V��P�+tH�#���<�e���:�mU>*�Q���VW��ZbP��i�r�F�>���:e�Q5͗Mmn�ۏL=����Ң���0�m`?��|�;H"��q��!;�g.�<�Z��O!g��=�>½�E=�'R�l2���TSF�RY��Y�˿l3�S,S���2蕏�RWѴ�x�X�'�'� ���.F���[l�q�`�*��Ʒ��g����G��E�.���u�B��5[�h�Zk =8��M���Ժ��<��z��wi�!�y�o/}�\��3-Y�𤬦�o�0�bu�J�.���5�\���7J�E��u{���l|��kR3��<?8����̍L�R��\z��(����s�+9��DRU�� ��]�G�$�0|pu$�c(HB�d����ر5$�����ƭ�7����c��uy�A��$j�<���5M�C�ۀ�K<�[�(�Ƌ�nz�GUz���m�q�с��(g*�Z5��H�����Y��.��@R���j4�(�ˬ�"��L7
Tq� � ��WR��/F��Ua�X8��.[�=f�12����SC����B��{��w2R�a����S%�v�e����9f"׉=�<�/f�ۖ{�8�ΰ_��*|�M_X�d[w��zu�"���ߺ8GC�"�V��'j ��?%�U��������4"5(A��x�hO���WR�S���\L�I�v�M���:G	2Tig*��<�s�MLik�[W�� ah�y���Gg�x�B����e�s�6r3f�K�1�V (�'���60�t��~t��H�nJ۾�}&�}��8�/3|�KԻ#J� ��ְ�ʕ���S$�G��/��|đ�f�8�J_�V��#�h1��E�"@6��fl��5.����mo���l0ޞ��5+������T�h>���UFB���IJg�x��ZB���io�3���J�n0u��k]Az����ef!�,.�D�g��.>^߮��j1V�ն���m�w��I�1�m<y��"��<y���!%��:Yb��OQD�t����������20L� c�ͻн:�}� n���D*
��X��W��`}�3_�����\�#T�f�3���[�"Y��B7o�!6V�@~�d��K��z0�F����ؙ0�h!�y�\M��}bC;��n��Nt�B�(���������:��UK`I'�`r����2RnW��'=侲�l���a�c�'�ֶ�H�R�[]��%ƿ��4z�Hf�_]�5�؄��4 O�_p[F+O�M4�<u��1�T0��H�m���S��K�}�_9C�+�∣.�=�F�tޖ0i�Ԗ����.F�D��Ps�U�0�e-�������?����@����^N�9���~<���Ż�+�^���U�ĩ}H��~��j>.k�/u��>Ȧ]>�żle��Ե,�����ݡgM@]*����Mϛ��QT��0�h��	+zϕ,z��f�ِ#IȈM�97�N5aH��w���}�z�R-q�J�����Un���o���0Ps�T3���)2�էr���cG�q4�qY���H��Xb>�)���.1%┿��|�,����tJWv��7hhn�0��r�T܍�x��jUX�`��=�U8��j�*`���&&ݤ��lW ?z5ѹ=_���X���Ao4߭�LRkE��S��",�*�ZMn���?g���fy���&�N�n��#�E"VYx��`e�a���i5�oF}(_�=Y���&��IФ�0�p�	�έ�u��6���Ӗ�T���<�ځ�s���:����7��}&�'g(��C&�UEHb>�R��ύ�)��HY�_K%\��>�s�`�fG�F�� �!���I8b�&�y&ſc�N�@Mܰ��2�M1l��������}
�J��2o�&<8]���bY�G,R��=Fr.{��_�ĻYK�r#����SP�Џ:isޔI��y$Ʒ�)�k+�gF�";��hȪ
(��[0�O�E�d5��h^�)���r���4��tzٮ*�8�gj0��"�T�W|)���Q0����'�*M��4�$'���c���(����n}���y3�f�� �)iJ��E�+u�(mD>�z�97Y�*m��wЩO9���(F�P�f�[?�������/E��a1ڹ3Jp�ɧҦ�~���^0V�bEK?؟�4����f�"lڦ�W`��O������%�������l�ǏifB�%0R;���l�U�8��NF�Ҿ:��s�=�I���}�Ck�!s�N��:Y�yw	��x�����|�l!�7'�0_"�B�� �T�v���C�hA_� ���W�˓��!� �՗��]'萅) ��_z	 ��Fڑ2ƹ�5���M~�q	BMH�;c({��YE~��uOp=B���z *{3k]�^�a�Ej����8K��\���q�߿M�y,ԁ���y��)�S�g�)N�*����]�a�|7�{���t ����,����ZϷ��	3'���8�l|1��he �'��>���Ҿ	.���O@�?>Ω���'H���4���
�\tN�ѡI�$:��tYj��~NJ=�
���K�a�Ԡ�,u+P��ߙ�1�\�P�I>���Ol�.,�1�޿d��Y����:�������-��I��z�� >��JQ������"��l����@���:H�7
�1���GO\3��{s�p߲�j�Ǩ�qAL�7�p.�u_�4z�N8j�!}���3�T>
\d
�
O�ι���5%E8Z'�{�ϖ�f��A�[a���׸_<8�O�)��&�M@�`����+�s#ޜ�d��FV$��+�������o� �OL�fXn?tRy`���y^�3��+�^���`-��to���QG����Qc�r�q����%�=��K,�ֱO]R䰤�Y�S���Xez���u��{������z�b���'�9��"���3v�d���LG9�-w�L"Қ��YXֈEPd��.��j����=������K��H��(��w�kIͤ���Ĝ�z1�]�ܦq��s�Y�A���m���M칩�g0�ɹ�tyOO�k�۳n�^A�~�Ƅ��fg�h4��p�V��x)�bI�+A7QE���;���X�WPIB2�(�r��0 �x�yC�k8��&|˄���rf��Z���;��u��s��gw_��>t\'08a�ָ��u��zC�P{�O��>16\Թ�i)�}L���&���>�����p*�{�6=�tjvf��q�`��]���4�)��i�l��DxԐ���*,�с��3?�n+.����ca�j��'�#�Ki(Z�!oU��B~���8C���>�QSfmNy^b�[�Ck��c/�����Q�%	�6@g�>��`3��*�2 c�����h�j��Q�W��df����ű3j
�����Ӣf���gJ���'�:�V&�d�Pؒ97�2�W�ٽpG�]��Wu�� �c���@����e�����f,���x���_�
y�:1�7 b��P��<���q�ȐU)�u9� 5�9���8;�_F>C�nA�g|�ӄz\z1^�禷�U'w��b�xz���}K��l���] �#��i�Q1�v8%��9���!ӟ��2��XqRi^�/�������Q$ۧ垱u�% 7;��b��/4�[ш}
��6�3�p��|�~��~3]ȧ7a��xvI���d"p��� 0Hݫh�È2t�v�ib��5]�.-&��ҙa��i~�� ��l���"�"�#�]z0���l��
��@�Ƀ/;��K]�{�0~a����bn�&jh��)��]>�*<�ӄml��5E�p�H�����[`^���c	>�w�+�_O�Ͳ LQ3$#�h��}���W�?��*�pbTxݷJk\KO�L���u���FT<��ΘQe�w 1H��wP�C�.�|S(��{��|����U�\r^ߥ+��̞�>��dE��j�R����_���[���\����A�f�(�5[�m+��	�UQ��_(^�W��� VxD�J�I�Р��S���⅝�@0�:�vY�C��� ��q4!���14�b����K2��y��zF25�/|�Q�(�rF��y�9����Zv銾Ǜv=�}��@h�s��oFL��UL�l��gh���Q��o�0�|:��s�R6�͹7#"1}u�W2�A�e���P�
��2�"=6q�,|���W���Mg�y�>���罜T�d�ng�aݥ��a&@b`�+ ����A��5^2�r�Ħ��Ս��������ೋ���8�;^�U�/�	��W�����1�'{^ͤ�r
fI2�8�)s#&�REl3O���LJ?=G�,��C�D�C�ڈ���'Bմ ���%XSD�[����db��bƁ�����]z����X�W��z?�i��;�P��I�6KN����ky��
S>Z����B�f��׷���"i��r�^9�-̼L|b�$m�}���4���)���VI-錁�N% �-�j�� �^pr9�!�Ɍ̋BQ�ϗ8��b�/����U��Bk�	�_4���̷�} c�Y��Kj��t꽀�:y f��{ٛ�-�g����A��)�؀\q��ϐd�o��z�o-��F�!6�/A�#r� �Ը6~AZU���$�i~<���Mr����`�hRC��1#�/�|>�����d�a��c��x�JJv���j�"<��u �݅}v|�T�0�z4���h*R��G�JWФC�C������ �!�0!t2&3c�d���&M	�?�a��o�!���7�ǵ}pX�%HC	��$�W�'H�c�p���/3�\��T�,�z�u���H�j,�S&��~VxJ�L�X������ߏ���Hl#.��~��^W����;S��	���'���f	>�a��]��9����>I��v�W�4IIgԥ�X,o>	,[������w"�\�v�E��A�)DMO?�8I�L�B�QU_ �@K;�Q&ȴ��)�9:e	��\�)��e������n!��8�ۦ�G+������7�e����b�i��"Y�i��� �u�stV����X����(�:o�7p�E�۲@���Txb6�^a� ����}܌��Eu�,�y0d�0H��Zdy�bLn��b */�M�K�B��fh��v_9�\����� ����pk[�.���	�=n�;;l��X����g�ѰpR*���Cb��}ݗ�>����u�ZsQ}�Gk�/.�o�g�)G~�|zISZ��\%��4�FӜv���+C��a��[�VC���&;9u���>����0�HG�A�7:�1R�[d��em�א���h�F��]�MƧ��S���T��$\|��"v�2�q�-���t�h��Ҍj�uv��w�Vć��VZ��R^�p3����1u�)�c	������!�����8�Z"�v�{�1:�)�76\V�U���z�v���JD�K�� F�v�|����Os�>������0N�_e;�����<@�6!(F�R�-��$Z��CH���g=e0g�q�F�m�鹧���/_]�mP�T��PF��]q_M�L��N���,�F8�E��D�I�A?+��i��.d����{�`�0Јb`BK�x��r>�0do�|S��E�O�*��秾@,�2D=�AF�:#%�'{�&
�7_�!$�t/k���N���a�3k:uܖ�|��^&Y�[��_��+rxFVm��J����k�BȎ	 �H����fx�o��6��ȏ�'��ѷ��0"�t�kw���=5�>&�갎�81 �c���	J����V@I��>���?����8�0�1�	s;rZ�g9�柙/���C���oW���# VY�UBd&����
б�4��B y�CC*Q"oHL6�S�fPG���P�¢�q��K�
7b"�rx�#vk�:�/��M��j�(��3%�j�4����C��Ř��@�D��q��
��b{đ~\�O�!���0𞍌�ϣ���J�e�~bY[�9��qƕ�b�[i�$�K���,�����N���l��>�m��<��4����}��m�Y�㣠�*oR��i=��Ǜ�' A-[��g��̡ZF�X<�=[���(�E�:�Y6�T4Dg�~����󏔱��LU�C�o��H�Z׎F��E�j�"q"�� y,[��?@(�d���I��%�-&�|�ZQĕJ�@�{���c�õ���	�������d���]�JհwI�TaS��ϳ3�Q��X;����
�)KE�5�B���aV->G����,<���n¿#���W�]�	%s0����lZ��Ͼu&0�һ�S|ݱ���:&p�?u�m@6��RA�^ɭ�&�i)�vy3%�@��q#j-|��Tl�(�'`�+8^4�,����|�Y�rvh�XTL�g���iy1���:�������e��z������̴�k�\���V���2,B~���/@�v�.�O�.������is��7"g�A���Ǧ���ȕ����~��֢��5��>"��$�~���Y�>Q��#�E�&�����%,tݰ��!�$|	Hyn�U���)L�����\�CX��-k���"ɰZz�2 ��g�1X��k�3V���.�&�����eɨSY�)��t*�NU��Ӧj9���P�
�|�?���R�n�I/H�������wf����&FB��ĺ�{�{G�Y�X�CgJs	�|i�E�Fv�3��A�N�7]7Uh�����L5<Kn�"��=9{#��.������б�敎�(���A ;��@s�U��>��O�F�w���ho�᛽����W�^���F=i沄h�}p�7y/\�б�[�7�V�_�%�5ܠd}]WaG��n�s��	�+�הu��H;�kIlMNq����T��#W\@K���f�{K�h�>8�a�\�`sM�28m"��zY~G�(B���\l�y$5!��J����ҁf��A�vd��ގ��I2����\.Uu�V��z�
�z�D���.u���*_<����6��Bv�8ܾ{�����U{y�|�"l�|[�
.k �	����淨˯�ZY�k�DΙ��i&X��X�C^��p�ތ�K�~���
�~�t}�wO��Z$�%���/�wN��@����2�������w�����&⻏���a������ᒒ��v��|�aju�'��3�=��<6��3t�P�ي�0�CW�<O�G+��CNq��~�@ I4�[#1嚰���kC����%��y�������;���� :*����Su ���V��7���q�V2�)k�V8��Ɍ���~�hw4�U������(�?3�'�
S�x}�tx&�I����v^ AGu��jH,�HU���=���A����D�/�?�B���SQ�<!��$�m���)ӟ_��� �[��?l���8�cǘ��w���L�a)�u`�wF��7AY��в*����䬇�^���jEZ߅\��Ъ>�
[���J4m��|�Jꨝ��bd��Yǡ�<R���O�	���naP`�oWI7�P'i]�\����x.?Ȫ�>�TE�C(H�:��Ey�y�S�%�l��L.R�/=m����@(�Z���T=���,wn���1a���\�DI�\-�����i�8��"���L�K��ğ�@h(��*V(g)�J�Pݵ�)����k�}u�ɻ_JT��r@J�Z��rxW��jAi��E�G׉UJA�X8���W���˕Y���������%�p��>����_5��-/Q�=)��9j~�^��(��F������6}<�5����Q~=�?�3��,�t�z�L�p(h)�GE�v�O�0ڜ�2�ͣ�l�e�N�Y�0��DUY7DB�hD�9�<���H�=��bh:���U1ׇ2�?����'��\�#BYP$vh3rB�7�}]PZ��2�DL���Fޜ��f��P뭒�K-M#
hU��F?�<͠�m;p�?w�Z�A�I+6�<���Y<�EIB��ܹ�K��X�����b"G�	w�ƪo+����C�`��� �o��y�]@yA��n���-1;��)�lwσ��5��V�+���mZ*�)���3#Ue�d�+K�׼WrR~�b@���`M��o'����s��)�V�v�.�3 uiԙS�T����Ȓ�hv�.群��A���mق{?��F~�MK^3�p�Ճ�ͅ��Dܕna�����;!8�4+B!��;�ؾ6$���R�	iи�ޖ���(�nB=�+<N`�?����o�X��E!�n�9�2�k�����re"	+�^�d��7��L����ʃ��1c�%Z1c�8�#�=<ߟSۭ Me��%��~���z��`�@,#nq��'�-���5N�p<�rt�zP8��13V�3�n�Y#G��a{����ؒ.I6�#d7�{w�������&���(�q�I�X���7&8j�ɟbQ?�HM�}-��@�2���,ؒ�x:�h���}N��R'�
��PU��?�9:�f8����1���"�{