��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�sg�ig �c��4��d�M����;��~"i���x��1�:��d��s�7U�S���\�\�,�+�� ��	�*y���3��u�Ӓ���y�3�!��j��m
W"{Lʔ̧"��ĕ��54��}ò�PG��ݝ�љFzҲD����rs��<�	��k����KMy&�w��kV���~��Ѿ�����s�B��ˑr����]�қ,��W6�����#�H튣�C�r�s�=.��:g�li�Y���*�[V<>�-�48��r���ka��ޥ�U{�[>��}�E�hK��������4	A
_m�՜^�ʲ��~P�'ۥ6N�� �]8M�.�2<Xr����!V�ci���eڗ����
�U��iwfz$�f1߁
8�}�[���j5��nHr�G�qW��v��)���	�u�CH���&n�ȃP9:�������!�����<��ʅtq���־܇�xCݍ�0V�׏�<(�Ω�O���@T$5�,�������6-�@,�`(�G[|�����7"c7�����pOK	K��n�2��b��{����+1�B]
Y�F�rB��M�N ��� �<�Vq�@��0{t�w���(j�������9a�5�Ky�gU兣O���]m\j��):�Z�q�[�~)�������c+�d��Lb }˄9�L�������ö�������G�-��Z6{��]؛ �3�ڕ&��u��mO�T%Jz�>�C���CO��1P��Ӵ�+yk�1�oueO¥�w�ѣp2L�ļ��A�% HV�p5^2x�O+2!~������Ē�=G9����ڛ�?R� F�}8�l�ny�r����Q}�
�f:7��z1�DP��~Q�;�7�C}�΅�`��}G�&�.&�$!X?~V+����er�R��Ri�>�Ǔ�ۂ�Q�4oNh�U,�D�I��+�|(r�=�8/?E���n.Ǳ���]���z$36�ܡ�1���
�3���zƩ<�Ө�_�dN�P�ʘ�?��%�,����C��5��8䌣8��=�g���j?�v�����/>�����rI��� K�S1?Zg#�����A�u���-c���7���v}��lV\�|ۗ�N�櫀��ȿ��3��1aL�t߄�u}:��j��	^`����U������v�]�:�}ׯ�p����tW w�+���K�K�&x��3W;�(�0����M��"���o|?�������}x��Zؓ��.�Aq�"��PQ��)f���<U�D�-w�ߟ�>���`U�AS���0V���� ,}]�9)\ȯ����M�eLr%!p��m|���R��O8�DL�|���L��w�4]t�4R�/��"�o
aI��P���2!���\�T�$��q:f����*�z����~ww�Rgz��'x���6cm�s��Y ]p�Y��ϗ,XQ�o6�>#ӳ����X�dIJYc\�����Ƀc�Ba{*�[mZ�7�j/6;*g��DM7WК���>R���p��j� up��+���2!��0x���Eͅ��:����5�.�/SZ��pLj�/�V۬^����u�������]F�naE�i��)tr�"eMӻ�Б�5�N8.�p�8�V�ԀG�Mm��Pƺ(I+-��kN�rJN���ӗ�ܸ�^N'o�cX��4̥O}�[��/�3KngOBJoxv��2�b�Wg���N�&"L���۬�̤f��ٰ��ࣺM�F���'�uE�~�b9cI:��r���)~6��vk5Lc�*�=&��Ǒ���_N�����o&���A;\��T(����끛-���o�p6���@����y����M�xP���?�<g�p���؛��"���p�@���`Ҹ��Dc�U���l�c��^�)�;?�8�v�Ί���w�#��t�ʙ���v8��q��E�5�my���6�H�Ӛ(��D�%�-��e"Y���������������P�RG���v,�,�Ԗs�W�7v�9#hA����-���(?�<���E2�B�2�����h��.�wB�Ĭ�/�$��w��Qϰ9 5LO�;�hV������tq�����L>�[M�
a�E��ppA.�#K����0�Kz�����P��l�R�y��E6b-0�I�M��Hdf�;�d���9�IO?Z�sj�ϯ��{�{H��q�U�o��ǯ+0��:t��)$��a�o7�Y8��	I�}����6;�9�@���!}`����g]��߮�ӯV�����U�QPl>�U�.���0�ӫ�#�Ā�M�a[A�"3��M1v�V-茗���g'-
m�����Y[ �w>2q!Q���"��0�S��L)�e9Z4����cw�8�T�^]��/%kh]6�5���G��7i��w�G=�5�$�Q�q���c����<A�к�����Ԗ���٩E�$�_e�{C\,�I��o_(������6 s�]��� ���W���%Y�~�Db>��YmX�uEU�`�1!bz+�p�SՒ�Z���t*� �{5\��Vr/+�����%����wj̳"��]���'v.L�#D~��l=��:i!熥�Ķ[�E�DN{DR�2����]�URo�xw>����3�@-��S�+��x�T�A���]��܌�M_&�A��J��8R"�0*���"���`������2�,��L=~�_:�щ���E4�ա��j휨��*C��xY��3�дae	@�H��I՗��'�JR��j��0�	�K�{��5c1e�	V	J��^8�0H�!Y�^5�;�̟Oel��8���{�ԕ`qaeY#��Lu���<b9������/����
����ȱ$�m1����ȋ���x�ށ��$�bG��zD�j�m�:�������`�x�����(�G�=��_F|��n�����俙I[.09a�O�z�R�p��:��H���,��-�(����W��\x���3����+k\��.�I�BA��u��Q0���\�{ϼ4�.�����aW��:n*]�jŧ�m�R�&��z����DWl��mQ�m׋̻�x�-�](1� f�#Tj0����]�qG�k�4x��:â�Pɜ�ep��.�;��/�=~�`d�#P�_TP�v]��Q�DN}qIS�|)8��������q���Z��