��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�X�C�[��"s�و����E��d Q��Ϝ�a�6+_�BC���~�;16F眵��bW.[�֤��%5�yY�v�U��/�h�*����m�0�5{Bǜ=��f�����~��2۟Yy�[�eYܕ��_�M�`�SAxiX�l�7Ʊb��{�θ��yk��X��d�4�t�"�HF�I5��Y�M���,�K���.��|��Q��b���zx��\��$r��R�2T�)q`)%�ŝ�2�w�u.��	�]w����t�JY����=c�ڨ�V9��B$���,&㭑h�T��"|ĒU�J�7І1*��E
qu���
8� ����t�7�g�ҵ��@X�:\^�mZaw�>�R�\�G�h�J9����U�?�c���br*��߹����S#��]Ѓ�X`꾼��1<�`�I��7��t%e�󻵸 >�η��3�X�y�O:���Vԅ�����Oq<Y\����W��kW13np��,��1��������O[��H%�0P��4Ӷ���Y�˛�S[aXЦ��ھ�U �����F����_b�	�EA�W�}4e,7�$��/���:]Jα7�dP�,�Z y+�HUs��J3'�T�FM�J�=�cs�
�α�U3�7����4�����v�-S�x�f�f@�M�S{�B�2�`��|b� I���p_���	���6ps8��s�8{���=R�q6'"c!铊�(|?Q����?�A�̄c�B(�J6�,�����b�w��3�+���yA��^�����G�����Kf]��������s����=lji�b	c��q��!8�C����h#z��k�
;�� �Z��iU�$�q�i��a^�ҡ3���09HV��ijt��i�\�W9<Q
g��79�X�n��+�kZ�c��IP/�?�.�-���'��Gd���5_W�|`P��M(h�0�}�#=�.e
��&���}����|���Уק��w��ָ̊�Q�	�;�Ǆ���4o��|2S��W�Ķ;�uT�1��E��9-��c �z�Ph� ���8�o9��0�L��0;�kI+k@(3�w�7�b=E�%;ha�$Lt�N�����u<
����v8~�%杓��F���1�#<�-p�n.��6�=R�"��>S�фB�Y�N"�&�Z��f!D�?Sv7�J1�ZXHva�<��bC	�� �u��R�N�0����u���Q����d��]�t�pr��ؘ�z?��D���a�؃�E���6&���_�}=�
�k��pO��j���N�t�V35A˘PI:��5�v�A��G8�������	�<s�w�p&N�#e4h�j�{;�UqV]�F�	�ȣ*���::�@k��ṟ�1eE�ڙ9��������eb�\ի�^l%�!Z�`��Z�N�={99׳^���k��Q8LADvM��?�?�v'�1���9(G�&�;���[٤�C)�2ΐ��٬C�RN��%h����0RvR�jn>��4B���^�ӿfE.�zY@�4峘��J�p�w)?5�7�b��!�Z���RG"X4/�[_oCD��|xc��&k�d��5k������aƪ� VK�/���q�,cO�!��a�C@�����+�3'o:7z;�k� ���D*���7��W��0Is��4�xW��S ����`u��H�G��r�tg5|ɤ��@�~>�$�^����p���=���G���Hr5!c `��D�,�C���!B���̈́DZC�߃���XyC�"d�	7���㄂��JsA�ٙ����l�Koh|G�G�߅�P�2N����l���O���=����/�Z���
'����K� �tek�u�\��O�Cv�j�hY �����$���>�/�$��?��J�b�lg�udY����]=�)�	��Й�~�Ȳ��Dy�s���)����7�@1"�?�9�⨬�Е��%�5�F�)~U�렗��xl�(B�Mm��/<!t�-��Hx'mX�:(i���\�%y�����$o�q� Z��w<�Ն�:��Ps�z~��7k�^kQ�´� 4��,�XE2} ��m{y�������U����&~3W�~��H���"�2�i_c���t<�P��I�`9�N�v!2Q��?Krs���C*�0�g��+��&� �U���-	r��#��ƙA��j�^%����44�.��]�_��̈́Z]:���U-�"�|�J:�`���7��9]OR�����_N�^�˟o��a<L쓣��w�2���b˸� ǈx�O��̾a�L?���/-7���u	n��9�	�J�yq���>��x_"��_��ͨ��R�(Ut�]HO���s�u��C1���ȞQ
)'#O0����!�H�>`l.U�'�ē�.���6��7C��V�s}�-�C��ܷo��Å���D�a��@W��ߖ�b��M�
�G&�v��`�������@��	�����0ԩ��cV�{��֪�����֪;u������;�"������"S���#f�~N�^��,��٫��\�$����wr�V;�٪VBf86e�"�����^Cv�o�f�)�����ppOu���N��b^�]H]^���C�;�"#Y����l�e�Cl�K�8�W�,�.t��ǁ��[[�O�L����/e� �{5X"��=�U����O��}��4j�_���*KL�GJ]����djPTƀU�k�O���1��� L��kv;���k����N:B���$�0�n�"�<��^����[����#2p�J�&��_m�)���")��7Dfr�,$F��р+��{���
z}�ܿI�+~��G㑆m�S,�#���(du`�{)����K�����`"�'�/�����xЎ���s��a$�Z��"-n7ֈ�a�.p�`�����1ڮ�ܟ�ho���A[��`L���uП	�f�����sko��H�J��{2T�t�	��}���l���{n(��V!�\���s��h�;ܢ�d^5�{��bZ��! �k-�X�~���r�����i,;�|�e��_e�+2I�,�T;����od��hr$4�N	�b���rw �.�n��Z8��T`l�`�R���-�ܺ�_G�ۀ�����HDe_������q��=־᪴	��) ��o�z0���5�ߟ��/D��:T�Ee-�r"�H�-(&h��DR�@~"�{�#��~i	�T�|�����)Į�Ҋ[z��Qh���ʯ��r��`Ѧ��E����`,&[U�C��S�sxH-O