��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�7ټm�lQ�חY���Q��3���Ss��t3�ɫ��zzm-!��#^�g{����Q�LC�k#��q����
w�i���]�k����X��Q#���U�[��åV�C�E[̘�� 
ݼ���T�.1Ҩ;�]��`�Y
��B�b���ۣ�h�ƣY­,��M$��sŷHٛ��r���cJԬ.��
ڸԋ��v&��z.㍐��L�H9�r�!�� @㢎!��
�f��ڪ-�!�����D���M�L���*�,��VA��(�k�@ijY$*�g����J��c�щ����2��qr;=y��:�)�`#Zߊz��8ʨ�*c���[����1Ɓe�L��u���˾������]��-z؎�b�э�4�|O,X��k��_�FB��8wJ6����}c,�?��MmӃ��V��0�O$�@��/	���m͞�T��������H|O�(����K?W���k���ޓ�s�Z�.��T*���WK���T�ƙ��L?�t2!�g�O:�`����^;̤:��8�zɵ�H!�̿��;^�h.���eu.A�R�|�Z�)⩢%F���R�*#PJ�|n���H��|D���6�֪W��W?����ªr;���]�DJ��ER��V��8�	������܇TJ	��lR��8@��gE#����*��^ ���UV�P5�7��$0����g]>�MF��쭙�	���O��D��θ���4�`� = eey>�gY����`EJ�u��7�x6�z�6���sxԶ/�D�X����&L	k9 �QȰ5L�i��#�Z����`a��� ���cΜHh,&�7�&�	���\��Z!�@���B�i��)�D�d�伐���I"A���n&�%��Z��ڭ��+ܲ��3��)�X�[��D5��*C�:���S����/��'/�7��B�br�5O��HЅk��X⎞K�(���}϶��p�|'aO��
EKmw�R����5��\ef�ھy�����3|�b+a�Skt�:[�S*�v�=�鄩��w	lұ���tu�$'VZ�T ?�-϶e����?P>�,<�����M�=%CN�,���J�V�B���Y�i֧�2r4�̒�����N2:#�3����:�P��[�g1�n�]U��fe�n���zs-�K[�/�����������zgb�3�n�<�4��ٞ_��a�jEQ׾�&��0�(b������1�����z"mτ�_KDwW�i`���f*��A������|��(ہ�42qq�͊UE� ���܌���[�Q���x�ֲ���T��s��x�b?V�x��z�HO���_r��Pj��\���i\\G�1���)<�{���=5����@�w���lO�iBv�&Ϭ�D����-����~z�z�!*�^4]��lC�U<�]KB�0��n2�C:j쫎��2�1u��7̘Ya��� 6��n�q	����Rx��D)\ϲ)��5$����<ˁ:;�� g���u8	�&��x��x�q� v0��;�AFU�Q8���MG���W1�fu�`�|�NJ�I��2���|���)��Y�����Z���_�Nl���>��9j�=��5�����mhʵ��qY3?��7͑��ķ�.��0�W|O����t���P{�&)�{��N�ϋ	���~��f.!�;����+�u�Z�[q�~����/�/j8��xwe��y���e��ҋ��<��7��J����mm^����5���CZ�����cǘ6	d���m@�M�b��Nټ镪����0�]5��?Zh�w��� �+�;�C��$� "�t`t��^�9�lƸl��,(kAI�� ��y���� �\ϯxY�4+��?GHiO��G �
����j
�%���=m���2���ni��̲]%h����ʸ���P�����l�,�Qvj�AQ�C��)�x��QEKc�Æ�m��i��PY�4��A����/���~a]��3T{�y�h�+a�ZZx(�f�H0��$���.f��1�UZՌ������8o6�t���~�ʸn�e �)��7x�T�D���Λ�׀d���F@ŸC�C�|X��&�֜�<	�ƪK����E@u�)Vl�WI�*媝jF�(��6�ֆ�$��fH��;�-�|nE�c�VЈȱ�y���|j�JO�q���_��ZX{��5NSQ�V���p���[�AV�r�g!��	j0�Vȭ7�I�\����Ȁ���*�xNnP����o)�Df2�h��/RF��
��e����~)=kX����!L��_�J�wA�J�W�륵jir���P<�T�#�9����ET�\Ppq*"yF)Ur'�دq����~7<�,6m�]�d��4)�:V�B`scMY�������t��<�i�)h}�E���VWi^���,�(d������s�����lS�v4>������`D>#���r?k�����Y$�H��r&Ƃ���9�;��L7B ���w�ci�6�����,�7Rp�֡ŗ�/��gR�������F�p|Nl�����y�v:
����$�ল�KY��\��Bcqc�=��r�ݞ��"�\v�C��DѪ�u|��A �^$ل��>y��)8�u��?�'�/��_���B��E)������'��줹w2��ˌ�\���J�u��!�`׌	���K`#���fq��gN��R�"�v�_������k@�7D��d�Rܖ̙4�PLs����z쭧q�**��o�^�;�	��]oXWK�1�Ŏ$��{���eģ�=y���'r��	s� ��訐��y�ƗC-4���fZ㯊�{!�4�~�c��E�q|u��/����I�2Q��T���y}iM�5Q��´�N����go-�23eȻ