��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��&�27	��"x�dA�G����87�p��� �&�ۀ�!v�#�_h[T@�j�DwҶ���k^�.��ܕޠ��_i���?��B�Q?�q#jϪF��n�u�?���L	��%�г��ӎu���QS9�Hmw���9�������1oH�M����4�z0��+|PB��S��W�xJ!-�4,!�M���3�M|[����h��B8���U�T�2:�v?O	?zCv�����I71_;�8 Z�~M���gy~؏w�5�2Fi��ϵd?�71��{�x�2��;j����69���/�⍙�^����
�ˋ���2�j��B���0�kˡz��@��9gW����CX��C�Ʈ"k���b�!����"�7��t)`�����'. ���J ���>��qvzã����L:7��(��A"_U��MQ�}�W�9���/�	J����i��|l�%L ���]�4�g�z����k[=Zi��a/�����{�?��m)mo	��+��eW$HJ�i��DApׂ��}���Cި2��O��ٻ��S�0����W��/�03j�W-�I�hEή��E���a�|x�О/,��iS�?�����1|�z�ۥ�QqM��X(���� }:�Ao�)R�K�lo���[!�do�����Ut>���D =�9�4��������I R�pr��}��C89*���a+��E����#	+J)��*�"Q�e��	�H�"xSO;E�Ј}C'� ��v'@^��4ɰjihtP_���s)Z�FN���	�-}��R�Cpě�����`�N7�vg
�M�o�^(�ش��H����n���j��\ ���a�2q��� @H6^�jJ�y}\�r=^������!�����4����2�1E���m}�K5��Ym��C���o�B�_l-��y��TSt�:���#��[)U��Ȟ�E�����3�<�rj����w�5GH]"ul5Ŗ�b󸯈�9�ʮ,XRA��N��|h*�b�[o�.�z�Mq��BJn��Ś�sT��ؽ�nѹ���t�&�D��bS�&���g<%��!���[��ay��\O�'b ������1���]�n�P��עV@	|�+}Y��t���J�������V*���q�n�h@��&�m�+>C#��*|dP�x���3�T���X�o�����e	�\�J��w��9���t���i�>������'���I��K�k霸ʯ�4����u�ܷ� w�:V����P��l
���D/��+�$��0���Lgqm�L�)������G������0]{*,��Nu�R��6Զ�Ҵj�Q����	no���~]kua3(�2W�5e`ov�2�� 6*��/-�+�,��t'T������!C�}����*����_N��Ǡ��GV�ɬ��±$��L8ҩJ��)J&<}:�Ja����wP˰����Nl�I�Lp�9Z�>��P�vyx��@U�p�\�;��N{�6�cn�'N+��fh���]����Y�ӌ���vD�a�b��F���3��B�[�+F��m�$Y������;=)*E�f�����.d�GP:�5�oqk�ؼ �E��b���ϴ�AF<���S�e�^Ȉ��ͻ%�$��'���{a޷4t�;;r�R��'��+*�iF���~��_�Z��Y�"���֩%}"Ri���Z�i����a��MX��!
=e�v�_����G�l�n�<���oL���E�������{!��T��E��2)���q��r#�Ǒ�)�f3��)3�Ꮸ7��}�{���!V���A�s�T�G�8g���^m���G~&IK���G�T�W3�Z�q!.�O5}a\n�6i�nn�~R:��]�n\d��|�����E��u'��{�nE�����$�NŎ�Ty�����f�ީ|(�.r�w�t��EY�槳Xבq�J:����G�.�qx��zǨ wQ�D��ӓ���O� ��/u��"�ؚi�����A3�5�nTGI+<�4!�K�D�\�Vx��n��Q�yM�+�h}���Aw2J���W6���ۚgl��' �1���*3��8�&-�ˆt��Ħ1�ɘ�S��3;���A֙o�56]x%���ݩ��Z��L�������W���Ĝwh
�fB��%$Ɖ,���T�V�>��S�F�$��Ӫs;���3X��N%d_geݨ����N�R���df���ɠ:�q%����bu��]��C�B����eߒU���2�`���ްԊ^�s�aD�7A'�j3n�b�\2��j�'�|�zó����['����jz�]�U2�k��8"���j^wNVdc+f��JA2i!�1�����R��o���-�/�Gi=��N��O	��9D�V����a/�Qz
�&��:z(�3z�ٰ�I�q��S+ak�-����,58�Pj^�P�P��*S����y(1|{QB���>\�M|�`���mN"�����߇���[�Q��4$�P�sI+�d����$��*��u�A3i������o� %��8WʐB���{~PI���[�UA��WM�H޿Ї��pZ��v9��1\�zFl�f�C���e#X�ML����#�o��%��o����m�P�՘}�Q�l7�6t������<b�cs�O�p�|�<�n�Չ����\/�^�_O]g*��ó��M����4_^ɶ
�n�v��l���Zn}v���[�#��j`/��JoR �b"�P�ƓM��<7�W��u��|3¦��׈�Um.�9�1Q��OfG�+�{r��^5!;���6\2]B?&�ڗ���Ʌ�������S��lԩtK���B����g�\A��3����9������%��Sׁs��T�nA�=�;4z����(����fSN<�Җ̭"Д�+��]�^��2Û�����c��W� :�Ept0�оٔô�Ѓ@�d��k�y��D�^�ؒk�5�;l'�pMW��������l�.�� MX���g!��d@�c��J����Sm���NYYK�Q;Z],&L�Sr����Şs$��p��m�Όd^����7W\b��3���>�Rϟ"}��	s�TM��(�R��b�7���,Q z��Hwf�j6��s��H:R�E77�IC�prn��a��ޢr��m�H?e*�~��?X�
���ui�z�f�����q���K����M�tMCXD�ߖ�ػ=
���U5W�v�}�'�|* x�>Le�~G���04�d���cX��qCrE$��I�h �w.ެ���}p��{<�>�]�/�����4���̲�|W�O�7GN�&���0*|�&`
قG�|��~��Jz�JU��W�:ģ�!Gu�0<~9y�^[�iװ&�z�w�1�V���Hq�u���I@�k=�t3������r��Rг���Ȁ�{~�MġN�]�U`��^>�@�2P>�gr���0q��3����ʑ/`I�Q��.����a�ڑT&���d��8&z|HbJ��C�t�8]�	���0;k�u�`�x�텃��c��y����S�ӊd揪��F�l��2���q���笎����&ஞ+�i��*~%;$ߦc�3��G	Z4������	M0M,�&��U�#�WA�̋���c��A��/i��:i�9;gD�5&M���ǽ�ǈ]KG&���W�Cв5;FVJe��']���~qeȕ�i�n@�݆�)�3�w�O��ہpu�o�4���>-�ܓ�3��`R=����/I��~���G��-,z�^�9�8���y���մ��T��kA��6�՗ɨ
�p���ҩ�2�%eO����]N;e��-�^���ρ�<u�%�D^S ���Ђ@�8]��4���|�,����T���S9kX-��k澛������K���3��n�����ma�*��}��qS�lmxu�������W<�X������+���I�u&��� ��%F�iH�)/Q���37)�yq�2`���_q���nB�K:}�ב��o��R*��r!Vz�N�w�O�A!i�����.Ǻ��̕�+A��l�$���]�q��E&�4ټ��H�_��L�n�n�1��;P�^�.�_��ȲgڼH>(�Ǽ�۞˯��)7M̖�^����(���U���
�V�G*��~�����n.�j�`��$g�b��}��nU�o�@�(�'�}0	Yٗ��(��a~��H��7�z��gjNE9�7/��s�W��i��FV"tX^}���%ef�nj�*��zɃ�o�8O	���i�or�s�����I;.u?!��V9������#��1��*^_Q�$ZYץaf�x�3j$}����PR0jE�?� X��v�.�t&5�J��i"K�5�3۷�Tg���]��ݔ�hщ(P%w��L/�nYj״AfW�6���X�eg%,"���._��B�Y�K��k��,y�Q��|Y�YYֈeT2�
X��lY9Zc���k��a�2.�~��M �Ȝ�|!�������jA
���Z�H�#��U��{z�m����G�g���Ÿ�-�
����i�����D� ��9��Q���Se`~|_�����).c[9k��Q�_Л��<�dӼ� ��r/�A�xH�&�e��4u��X�eemƢ]lSp�!c���[P���Ʉ�@��e��-�I7��8�)�l7�n$�=+K���Y�KǜHF��،�5�gI�*�1�
�J�(>M)"�]U��S�L��	�0����Z�Թɑ�&��U�l�y�^b���9�$[��!����lB@zgA�(])TW��;��vG�ÙYb��۳R�u��EJ�#�b�Y��sXS���_�o��E8~!U�d���-_�m��(���Nm8�z�iiJ���nx��䶉�8���͸>�7׻@��㐄~�i�������b���odf�Xf8K�.�����E2Z��@�(�<��i�e��U��˧ph�Z����7%W	�3]	�9	@f@����M�ISM\�7��2�A�J*	���S�apۥy8��*�)��<k���%N�?[��ߥc�a�3��v�%���1��l�pM���Oz�cFA`\���<G�ÉZ���C!�0�`�J���X�b�\��&�N���ד=��_�@MS<v�;��z�!"r��&e�"0�ݪ+�!�Z���]`��[�y����|����m�~����<iI��W�E�i�[�e�(A�OƯ��#ͮg[ZI2j�M�r���$b�k�_c_!VV�eD8Q���ǑV��l�k���f�GQ2]�Ot��j����yy�����'��4�&�-!e"�G���!�EE�!�ڔXw�F�v��/�4�	c����j��^�Ux}�Q�2�;�yE�0xuz\�A�R�:���b�q-x��#0��\'y,'RQQ���?h2�_v�Jk�V0��Lquث��.w�u5TF��U�ۭb����w�(7��d���4�4��9��4�����|��^ߜ1��#?�Q�[�uoM�Ȱ��a��:�Ţ���<Y�8�� ,[�lˏo�u��D�v7�z,��[�# k�f��\��_�k}yu��L���I�b8����z��E{� �w�n�o���"W�˷{~���˛�`2X\��V�b1TT�>j�TSO��/�sռ�+�B=6������4�,�(��:�X��m�5������r¦�A˭s�b� �����_0����<��ފS��Qm%+�$SC/���ou��DHN������A�k�N��
�9`¶��X�kͭ兯1�0m�½�e�t޽Gk��S�"��K��w�b����7�8J��_d"9g���;����U��z{����´d��='LK]�{>�R2QN=�w\*�K�J�|K��A��Y!h�����h�N&��J�R�XKT����j`���H�7�ڀr*y�F48N�xa�����wDF�U��l��&����O�T�@����)X�i�T��te�Ƚ�M�ԵL��K���}ȥ��Me3���h9��Ap̾�-�� !Ѻr��3S����V���ay�mP�(��W��Jm�;Ŗ^���N"qU���d&<2�E�P]�r=�9\�cz��4*|�A1�9����J��[&�j����g����뿈��Ԅ'�^-�D�i���f�װ��Q�����>U�M�Bֿ
�q��e��˧�i?Ʈz4�t����{�W���h�c��.C�S���ӽ>k#�iY���O�K���Lۛ�Ƹ�fd��0x�ね���㿑O�`ű̘Ѿ��v`� jd��'���l�m�a��������?��[��\�kZ�l�͛ߨ��n14�I'�
�eg�,2�m@m���ڸ�zR/Pf`���N��؂���q�%�����
L����XV��8��3um�s�bM`��t>!��W�PЀw6�0�'�d<��r�)�`�A#�`Ѩo�p؏���3Íh��ϥ{iA��;��?R�{p?��.�ء�&������YΩ(��\b�!�tS�c�
��2)��dD��R�V%���P�%�i�������5H��͜�id�q�S�����2q&m,���U:�'[����7��ڸ쑮�u�\��և�i�C�9}�<�=�z!�n�u8SOr\??�]m1�[�2��8��\s�(qC+ ����[z��řJ1��]@E�79�2ჹ���1��h�OB�v��_�6����;]=�A����i�%��,�5�n�`(���0�&�Nfwwo4�s�{/��Lұ�Ÿ�[%��/�gѩ�B� ��:��K$�x�[yU��+��p_�#��v�Pt7� !Lk�~�,vx��M��L:��cAA��e�x10��ņ�n+�s�q&�6}r�S��"q�xt}(*�)zJ��� ���K�S4�x�z"��u"�SvT����%�_}}�Z������l�����NU��/gw�p"	O���m�P
_��f%�ˍ�q��͖��)k5�P��<��A�Jε;������]¥�ۑ���SJP�"&�7�����������a���E>T&a�������>w��}3�#D+y���C��*�y����d#�Q&ȼ+���2���+�T���ddrޞ���1���"�˨�H&$��ؓĚ2��A\R�ܢߖ��H7�7`Y�E�jFx͡�������04#q"�I,ES�o�y�<:�P�lP-�K(5��Xy� �o�[ϲG�4J_����[����j*��|��oŗ\���3��.�ӈ��и��`����y�g_3%�D�H��j��Z�Wޅtj�1a��b���Zϩ�wj�f�L����n���TF���؝9�n��?qq���_��duPv�S�ܔ����UoA���L�G7�E�Y��ȯPV��yh���N�:�(�m�T� ��+��Ss8�W�-?�5F�@%��4� �NO���;5����wk����������!<��cҷ�GNIC�ѿm類ɓ�ޜ�C]����m�;vf%zQY�Ak2��^�b
�t�=��U���8�<�:��ٜ4��T( �����m��PZRUoM>;�n�hkW��SKT_ Jt�l_�Z}ֿs�?�m4��mud��z�J@�}JlQ���!|��OVg�G�a��=���������O��(����Rf�;9��:8?�4~Œ�'5�x�P�=\�n�\5T�Y4q)XS�!�Ӳ�`S'��)`-Os�|�cS��:<4y� ��ʤS� �
ؔN �����Y��/���U�bL�����]i
��Ea���[G�ޫ/1�X�é���oև淓�	�R�OSَY�bv*�{رi����C0�p䊻ԝN8uڂ��;(T,�*p�F��
J�H8;o�E�m�5�nsSNYq/{]��UVa��%�GV�&B��P�tED��鐛K��y&�;b�ɲ���y�+!-?�Բ��Y�5�����IIo�ދ�c�֌B%�?x[rS����9���!���b�X����޸c���?����;����"�K4�ăAs@��{w^;.KE����|.�[)K3�Y�H����ɐ���4��A����^���Od�9�u�P�Ofw(�,���v�y��$���E�jaZ�����������r:ɠ!�����i��-
ÔHwUL�(zn���ĝ����TBߞ�pT�ϋy���kdj�zi����(�;�n���
��2-�� W��cy�-�G+�*��Ҥ�ݩVfd�ԩ��*��ٸ��)��Qۗ*6E:F=�ZNa���P ֟&&��̍'�q̠���lp-�E��-@R]���k�^��x�$|�+�J����a�\/Pt�s�j
�G�hi۠[L�s ����F%֣&�.��uC��'>��ꝥ�Ӽ	"Г�[��?ϰ��HDJ�,�Ҥh�nF�KT�|�f��x��~��եlpy�>��4����8)ǣA7QT�]�V�tX:Bn�/$F�F*� "PB�(3	���va�f7ss�Om5q�>����I�rL|"	in�@��)�z�4&kIV�ã�pQ��YUVy�q����s�:'7L�b��"����XZ������0PTђ�[�ڪ�7k�J�]*�)Ո�oO�e��2z�t���G��,D�t�[�3 �ÐA�	}��)�E&/řN"�(�y�Fx���S���3���i�0���5�ȉ�U��^.�))�J�ң;�v����O�]B)���؉���5G�B4�����{:�=8s�C�C<i�4[5���}����kӟ��_>(7\ R@���Pְ�H`з�?e����ɱ�^s�K{�k���=2�C>+y� X�d�����r����i6�-*�]"�
E�R�>�|�I��5#�;��ϝ�zg$b0u�4��j.� "��¸0S3��a�!�ć�"���7�(<�����H��6���>x��ɩ<Z��K�����a����v�`� �[�pԯ�Uj���p@�99r��j���=6zu!Tގ2�"k#ksv	Wʁ:��#-�հ�K�aPL��6y0�S�7%ˈQb�bI��I����Ü>[�]��E�BC{�r��H,�\�ԙ
�����U;!���QS�ev�ej4�Ј����P��⮀�}�͢*���V������/(?���Y51="B�{w��,�{ Ƈ�.�NAc�G4�]Y�3�n+ 뷶uzN�{`ǯ��u�F��	4�\���«��՘zJ�A}1%�h]�������NCM���������$Z91?�	���1gd�q;��jL;rP"��p*�lE����2\�RZ�5��ݶ~�N-+�3�e]��کh҉�����#C�wx�9["�C�n������#�~��	����}�"��R��G����8�e��"�BA���Q�y9��5r��~��]m�*G�u9 ��3��?�w�	�GM�I^��b,���n�V)�I�DY���ЃQ���|��SrB��d��j� ���,��\W%^Y-]�&��Bm-�f��8��--����-��Cz�$�Rz!B����äq0�
Sh�7a�
'�`���d�$� a8�N�8d��8�\�si6e�dkn�$R����P]�5h���`?jq���o7(d`�ի����ΎM*2�	�u��8�$q���j}>a+l"V˨�!a�r�6�*��{}��\p�xCh�7��9�W"@rν�z�є�*��?-�'���㌜�܄g�Z!���U���@��F�vt�:,�L�w�h��~�U����S�s�����ѱ��cA� 2�XUo���N��uo��4�>���L����~��^��]C�b�ߡ������&|N�b�@m"���m0�zr�O�bA#�>G{����a�`�6/�Ӭ��{hM�R�f@_��E$�8( �b/�T��mT���Vٕ,Sl�]R�ʇ��a-�b�@W(V���w���)Q�Y�Q�:�� �7߾V+;z�`�C�?��mYp>\�~��z���a���k�F�M�a������,�~�Yk��Tq�G����v ����ۋ��/C�� ��8$	���/۟�&:�R��{YP8���-S���@]�c.�W�?����ޯ��E�9��1�+������rr�7�-�Ǡ��ÛV��_�4��<�L�= :�~$q\�Á4�T�F����(��'�0��� PQ�%����*t
ޑ_m�^K�����Z8<��b�}��L�@�G���H�h�,hY�aM淶��8"�L��&X�J�Jk4E����yp? ��Pmx���>C$����
�@ [2Ƹ��k�Mó=$���PC2[���<,a��,�S���C8��R��{&o��v�����	��6Uc��5��ĵv���O����+�
 !��"a�;�P+g��hm�Mx��݃P�>�2��	�85	�b9h�ު3X�#�d�Fz"U�P���ݲ�݈_a^�UE ��t��(p&��-]��X���'N�.��������cG�	Dt�����j�MuL�/��e OZ� ��ׂ�����4=?�0����T��v���0w���CQ]+�G�l�`�j���M�o`�V������+��aZ�C"�>]���̛�1ff;��ĕb���_����1\m�*��ġߨ� 0�2�����M����tf%PL�Q��_뾠�g����	�c�<>&*���+�Ǘ���,k�Q��U�)ZxAB���ͺ)��ϱ�&ږt�U:���u�d3!ea�sP��36M2&[�������V�s����k���Be���\�Yt4�&���1<��u�L{4�vH�u�HA�s%%����0ٻ�~��Rѭ���7��u�