��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�
���B�+�����b�k�t<n��!_^|�0C{����+�f(���͋{���'�*�
��(�C��5���P-E2"*��t�[���E���E��dZ��J�pfq����@\�m��_�(�#x-�=?뜿�X�(�N���J
�\;&�;2"�%�ZV��,�؞n�V�h;&�j�!���X��i�bZ�l}M�&�l��۶�Aȣ �6u�0x�-�����I��a�>q@��l��;�y��s
�5vn�����)�IJ1Be�0�E��r��\���K�UH�ȫ��h\�y�J$�E��asI�n�0�0�X�� G�x��i���dڗ��Q1D�hV'��{	
�}�e)#Sг	�`p�O����s�\�5���?��۲i-`$G.*s}���~e�X2lF{V�ȇw�j��*����,�9-}���C�Mr���I�=|�{���|%��0�-m�o�~�=�)��1\=w ����Z	�qn�Npx>�V:V���g������'�&����ly�
/f�3�6�ܮ"3b8CXZKD�yOӈAi�AA.0K���%Ğ�����������T~�VqW]�hn�}�FC���)�A�ĝ̲�D��@۩$!3p�A��/���<��U�ǳ���������H�N����JvU�pu77�R��C�_�h��ڿ��/l���UͶ�>��2 Y�չ��ǜ��f�y��>⥋��1�3ט'��UbM n%�8����u=6��z\ʴb��H�*t*��=)���s�C�j�+q]�]�6/%�x�N~��c}`���z'�XV�C�	����;$�澊H�wi#2�o��0Li����2��B�m�7K*�z�%����0~~���:I�j�_l��*(��7��u�� v�Wv�A�Nw@�o�V��]����=�F_���w�g�G����,�lxd�v����p5D�^��;�1.;˫1(�����O�>%'�¸��1E��ꟴ������Ȍ�t���~��\b����{���~,zZ���-*�&��6���x�!�U�Wqe^��˺��7��t4X!���X�fG�:}|7�L��!�k����,޹;������x,�c��?g�%o�1A�zԢvu��AZ��_�m�8��R��DW�����-	-E�LHL&��'�x�:Ũ�Q�E��O|� 2�Iq9p��{���1ZB@[?�[}N����v��%g�=�������Y�ff���%;c�A\�V���2B�L���I�*���ͼv_��FE}J�5H�T���2�>8�q�hMr�Yoܺ1�����o⑘��t�B^H��U�����`� � �<_w�O���h4a'�|�܅���$��@*˜I8P�r�2�9�g{eh)����&o�.�/�����i�"���Ec�U�7�ȇ1jya�Yg���>)��q঩Ҁ��.7�`��.o�T�J��8����W\�V;�і؆���pG�^���R�M�O��)�����'C����y���h�Ѳ�sp[�[[�I�y�O[xC)Y���Bs7q�k�&g.(z;���>F����3X���gg�B*�����9�`׶}�P��>��g1�;ȍx��繡��k�"ږ/�~�4�!,̲c}�3`�e�7����fT�cӪ<ϰ%�����ϣ�5����Wu��� �6�9w�չ�+���;1���}�'�)�T��Dȁmu#��V&��_C*�V��N##fsaDH�����l�<�u 
yΡ>�ߝ*�	���1h�v�/4� poTH�RvvW�C�\��˫���_�c����Ԗ�E�%�R_�X�y���{���v��p�:��1�]~�����]~����m�!.�{赿wa�jo{yy�ԇ�V;_GHi�b�������M����y��B=%�����Y�t2�A@�9&��x��`@�&ɻc�������#����I���T04�huV�h�~�h�:jP���&��5���So�9wn��F�P��%k��Y� }Bɷ��
�*�}gYd�!A}���9*�Xn�DӉ�q��B�I!P�p�
��d}�s
�d4�F�2����c���\}���QZ���R��f��B!(1d���LW=��av y1,�2N@����3M�/��h���!��E�|8�M2M������S5���sHW��
&z'�	bQ/SI��X��cC�D�r
e�e�`-�J����g�K�E˶��c:����G��������G̭�%���p�����AB�kE(�+��T'dz��F0��]��Cr��� 6:d�t�@�6�R�(��,��/4�G�G��-��p=�|;��	�|�����t.K�&J�\@ f(����t&
&���C�)���F�VQPp��~J�����'�$;�®��9�8d	2�R� �\<A.��*��Pdh{,3�F���0���!��U��֟ ����"�US�{�O�j���U�*I���n����z�����+3
=��(T�8�8^��"3ʾ��!���Wo9�_�1�M����T�%�f׌�Qc��U�5���MdoX�\�?m��齽h���=���������	`����9B���E),���a��"�(M���?�Oi��X����}XX�+�C�
�3�[e�f����}���_����x�${]0�A�T���3.m�w��d�]!�"r�w��4�.M�޼���x�*��U"�6��Ld�@����3����'y��z�G�Ow�Z��sb�,m�3�o��PS�	��Ν0���)���TBq��Ʉ,cdp�oA
0�à�ٺ;s�9���[T:ֺ��ı����W{�?��O5�4�# -{}b���Tڎ	g���xI�k�-. #k O �	��P������pv"@��I٤������������ �Ҽ����G�Ͼ���T\��2�%��s��Q��]�^N�r�9��Ǩ��c�>|^	~(5[gQW�DM��>�	 q)�ش�;�Z.�Q�N;I�E�%
^��(����B ��s��KF!��3�Ѝ۴�s|��˪Ntvߖ���ac�hb���C��z�B�C��� �m������zI����6Ԉ	P�|��)�6d
�Gq���z(_����
��pf������2������G�����E5�n��Áw��K`�l���)�ba9َ��/֍m2��+�Q&/�op�Vw��鼌#�U\�dND͔i?}��k!p�}�0���5�̱d樔��uM�T�]���e �=���e�Y��Fb˾[��$�K��1���?�l�gDB�� ����l�˨J �gMN����%�w�y /�a��i1q��iZlr�9VF���K��T��ͩ���^��A2�	1��e>�!���%���f�co����fE�_$HNd~��o��&�Z�IH��5rd���$�k�د�b=�S%���^�u�Z�js1bk��ˮB7�e�m`�b���u\�)�M,�U&�PJ�
�v/=���^�a;Q�,�����̤����<����YH�s��A�̨���J�t;8�^�Y�U�� ��n���;&�v��d��K�vX��$)%{MXE;"~+U�{����
�� "�^�X+��@*LTq�ˁ�/q9h�8�/A�B���,���n���v�N3�zԸ�=�-�~�|~���u�S�;s�Ks�9�<�=��������VdsLt�Fo%��8[���j
2��S7q-��O�$�Vj�ržTG��c7%}�_��纄��ҙ5�1�43����'�w1r/�t�*�t�h���]�w�4 dv�%#�틀�KH1��'�H$A��� '����ݽR������/[r����%W&�<}�:=��<���Q�_H�zv�b��%?���,��畏��=Ȏ���1b,.L�i�8�k�N�j�kUL0:��d$�0���4�s�6���_Up27&=��?�|����-9�d�5c�S=;�lk� x�qG�V1 �4�:}��c�+�&["�@��mdWo���&?5s��9�w��a��;V�U�kw��vy8؀#<X��@�Ʋ.tD3W�2�`��)mj�a@�WT! ys����+*��y���+E1 iX�3���y[�t�$�S����ꭉjHL�r���˂�U������H#tW�g(/Fj���Y�*�o'WV���&��q�Y��f�G<1�����8q{E;(�@���+��p��=�� �1�T%\��ߴ"��H��c�B̢#���#���� �- ���7Ď��7�Q��5@%�Ee0�&����G���r7׮�w�ޫ�㤝O7�Mq?%����#���o]���ū�0�"�����(�SW��8�/��#�p�y��V p/C�{)��蚟U����ߙ�7�ݴZ��UM&e�$Ͱ�J�j�L'������WI�6��9=%[7�x����,ؒ�]d�㋊v����~RЏ��(#0���6��Oq�'<������[�CѬZ�W�@�%�y�7���ꇸ��R`��'L���i+��B�����t �cM!��5N��X>���$�[#Cp�1���w:��A7ap��,9:
~ޖC�:;�Ex��e	W��"O��2�O�[s��%�H��7Fɝ�� #��N��N�_�da�5jJV��D��_bԼ�"�(w�������nOrf�=%TUy.)w@��U������]�x�#8��^q�R'�7/�U��eLI��r(n�l~O|�̳�S3E,�	��ʋ��A=�|IQEM|��pƧ���R�Y�D`�B�?A��4����T�щ=N��L�jw��~k��/Ҟ�o��֨������<U�Hi<��^: �0�����7���*��/0XeL>9�X��GR5����]�J[��%Cᬩ		b��6�~��~	v�@)�Y���X��o�h)D��������Hm*(J�W2 �����
�'$���C���2:J>ȘT��hc �~rP���ºG�����a���	�ZU�HV��٠��P��BY�}*I���	/��z=?��@�>�"Ö{G����~7�}b]�ܹ�B��(yfiSaz�LY\�F,:q��aub���eٲ[%l�e�+<�-��I,��0۾3��K���sxy�k�����U�Tl ᩸�����0���ï�U�q.���{k)��S��A���K}�q{S�IͺQ�?�H����ڥ��Y�vw�P�!�8ۚ"W��Q��M�Î��F?"���/H�l�A�3�V*<��]065�|]m/��kZG�`"��`^g⬿&`"=�Co��D��;r��k�e�Ųb>d���|�+�&┺�el�gD(��(<1��'`<NR�����en](�<��Sz|9�ayb��i�%�Ҕ���_����h�J����QV�w����XUQ�iQ��:+�@?Ӆ���zW�{��}'�}��b��Cjc72�3G�r1"~uWx-R��Y���qo�]P�ݓ�,n��
:���t�7XX���rz�� :���,�.VQ;���J����T��mG9�)3=�� ~aZ�DV�<W��i�������uf��[����6�]c���1���#1�&����r�rI�ʑ��=rft��Wd��W�MS��益	��!H v������yX��&�+ɶ���Zۮ�S+�q�/��Ta��}('�]1{zS%� �S�Q����Ls����J����ɸ"���9Zr��@�\j�u[�^��@�*��Q�$�Oe-},Uv�7 M������,=q���3�2�x���^��U>Gr�b�d*��A��$rU|徯�K6�ݝ��]��H�ּ`�*���s'\9�����J)*:Q�f��n���N�Po��X0;K8b��k�|��^M�ש�7M��O��v=��Y��
Tӄ�+�������d=���߸�.��!`ʿ�� �(,��.�th��Bc���  �� \�z�R�nCnl�I�����I�ʚ�vq��֋]��t��!�.w�L�l���1-C�m����.?F��4M��;c"'^��b�(Z���EB��&�\���Գ�$����Y�q��y��WW'�"O����~��j�\K�trc���,|z�4����)��v�$$�H
9��[��?�K<$�\��%�-�o�`��}�|�"X�\+�?�i�A�H��K��l�R�9�I��Y'ZT+sz����@d���:���	�X��uze�\M:�AM,}���7�������SO��tQ��9�*�վ;bwKN3f�j�����+��M��:��cN�=5T���Fn&��程���.��%�㊓�e�	�)�<�H��3����-�7&�BQ�놱�B+���������#���]��ݛ�:IX��_��i[��:���e���-��za�<��}�􋫝��)m&mv���*�3G��1�p:[�+�mR�Md`��e;3iLH��v�}�Ÿ�w�D �-e�]�Y��VJ��i�?]�_���9��Eڹb��Sđ�n��k� Ɉ�� ʒ�0	���=]��e��3S���ӝS�MGܖ�GMô�miog>�x8��0I	<KΈ%�2��_�s͉��	���#'��9��iݚe�mg6���ށ�#��(�� �qOq�+��)%�����/�~�p�-�y	`�ǆ��c�	�Uy����'��0|^�+����J�4���ږ[x4�ܮ��t�\�,':UO<�0Nh4:����7|>� F,����Ḹ��J�ķojnP\A�#0��H=��X�F^��m�43�[�w�" &�����MM��K�d�u�����J��ߏ���ʏU�`bY���,��H�B�2��T��#�)``N�1�XQ�͏�Ί�����;�$+�^IlxVĩ�$)š33䀄eИ-���@�;{��6rnV�Z�.&.��/^��Y�O-���N�l��>!b����.�ɿ�����j��͇r�u�UT��`qR^��� M�sW���sF��P����y���'��4j��Lo?�E6�(�����ķX�47[ZO��d�=a!�s	�C�\�(B�z�e��"�ʔ���-n��[���q��,\i��1�,i}�ceo`6�cG���Z�1�xkU�ŏd �R�́p�e��Bų�֬*F��c� ��>	�H�0�:Zp��aXQ��|҆?)}�����$nζ����U(V�|��tZ	�ma��;]��fÍ7.�Ig�ϕ���j���X}���2�q����;�۔�����0 ��rB)kn�",������Y�߾��?΁�u���Z�����[�e�ܓW�P��Ӑ�蛍��O��f . ]��-��:�ad��3���j���Z��-��%"./ZPeߏ*8
ċ`��󪎳)w��N�q��:��ٷ�bLL��Wqw&�!�/ת����3l�q�G���_�]Ko8�L�a��J�+e��>#�=�P���dx�'����������q���3�v�	�N}{%]R�}pF��RF�ʈ���������|��@��b���]�(J-�HR�7�M��t��L��F�F9�O�?*ev���'�L�����+/�ġ��:��jRx�$��Đ��GT	�����W����)R����ɛ�����wM��P.���t�3�����^��8�	E� ��^����e�Z&�?��2� z_0$ÿt3�&bҿ��L�&�+oK�[�w��V���Y?/�/��G�ˆ��
|��uh�
c���r��f�sم\�v��"�P��O��
�	��!Ih�o�ˍ��\%D����#9k���!c��de�#��?}���9W�g8�"6�H
��٬#�KPm�/�F�'�]s�����i|/P~������̧�0�rC������Vr\�%Q.)����4��Y�ȏ�J�ўe6�zAx��D�1�]}G3/�e�-��a���=�"�I��SJ�cz���y���α�l��ʕ�v��h����N���ߗ)$IL&�#�6@#��6߯vmN�e2���Cc�T�%ۘ8�z@�'�
����,�}��0���>�aDo�
��y���ƃ�i^KW��qḺ�� �}�&}o�Oq��@j�CDs�Y�iq@3��T�T��&hO7����Ge%63�)�=�{l�)���hFQ�F@��vf1��EA�,`�2�u�Қ���Цj4�0�p���k�Y	��_��q�5=ed���7K1� :�W41�ũ��q�؇����)��P��3���9�p�}�!�n���_�>X�6�:xQS+Qk��b�#����~��=����+ż���-ͧ���ÿ)%�Mr�_;����f

rk"�!W5<��x�Ǻ3@�4T-��ᡛB���m5D�e�0H�V� ����]l�"!�7O���7�6	?=��&��0׽ڠ˰~��!�k\ӻ;Q)��*�0b�]�h���^�c�i����~�a'O�;�����?:8���4a>�K�2��Q��:��{�<ݵ�����������Iҟ0��Oia���J���V�瑎+&�Et��-��t������ڌ���8�U����^8��!@��H�Y��ھ�7����Gu��#NC�!o����7��P�2�!Ct'=�~�1f��P�LCk���x����B�G�)]h����
a6)�.L���"$)�#����Q��C�����|o�}Z��Q;��?�˨�ky�7�=k2A�\�8d� � �UP�6ē�@g1z��g�۳b8���T��0�(h��c9jS��=�Ex����'|��*����:�6�J.�uEX�[���־@��'b_�;UC��o��8�I�����U��61�7�/�P�f �P��l�Z"2ȉ���~��q$;��xe��{����Z�*a�f�KUU�t��������4Dj�T�j��^b\���U�5���>ς� Ks�Tl�<fp�.�1-Tq�ĭ�,��!94#�e��D���'�^��5���8��	�w��(:)X,?~(��
�ߒ���W��̃�Ք��v
:��7~�K��4�ں9*r�?N j��3�rP��IN3���&t�T���c�����mJq����7t����%�	Jza�l0��Ayt�]l��P]���5
��֍�v| �&1J?�����^} �P$�M]xg=2p�3���`a�?-�7,c����2���0DE�-�1�l��#`:t����W�ך��l��`��y���������L����MU�|@IL'���m���xaI�3��̏*�e;�h��51��Ә�dej��+�7J{���l⒤��y�}<	Y�*H�"��^��,�'�^@����}~/y
b՘��%�4WM�0�%�(r�]2�;��0�yϤ�@�6�b����s�t�K�̴�_	�ȅ~1냗����3����j�_QA̓�v�ob�$�A/��s�kq�2*�cU�P 
��bB6�O���	�y�w�Q�U�_��%i�j�m�_��;{ҧ��Ơ�pfg���9v��H�2F<A�b��N�Az(��ޫt�?��qt�<��g�-<��H���
 N�U쑃�-?����woUU\N�.�I��Bpއ/���~ᷝ�>"��QD��􀋵V��WQ�e�� �~,Cs���*&��; U��Ht�8�o  �'�p|Z� ��in�)����B��xNOv��H�b��]�vh�s��,�N/���|���	�HT�)榫�Y�w����#�N����'}���BF��!S@ja#�R�K4�$����5Y#XOb(�5��p�7@�ٷ�ܷ�PC���_:6�<e(L���X!�rXh$�0�[)�ф�Sm���Zo����B����A*֔	�V~���`=�>��Z���p�ݨjO��_��{���>PjSj�t�S!���;c]�)WP���y��f��D��M���h��V���d�lg�|��Q��m�d}�۷�
�-��ß�t~�C���9������}���]��:��g��w'��)�,�m\L���D���KU����r4};0�C�~z����F�Fa4)&��M�*��_Iw>Sn=���XSn���F�57-�_�:�_����3�3���@���">ύ�x�)��PE�z� �'e�b��q�@*���qs*ˈ�n�x�c�ι��)ռ~@J����6�<��ϫ �`��N��j�)�p�Nd@&8J��^����� z�"OX'��9�J��@��z�5�VQ��o�Ip�I��v�θ�[(���+X/�4�\̬���!�ֆ��$N ox���'�Fԛ�ܦ�Kn����{�~g�qj���<�<8��=�F�on��!��Z�(I#W �f�0e��CT������5�C)�� 6R���QM6�ILp%
�?�h#�n��'P6
Y��|v؍-�i�t>�����*	�*t��CpΫ����}�r�'�B.��=��-H�!��k���k.�^�|%#�=�FӭJGpA2B�d��	��f({	�A�s�`X����vş���۔)X���}�Y�-�*���a�o�H'Ű�1��j���rlM�/�����܉}J4���d�q~(j<1v�@���w��f�0����������*��T����=WE@�򏽬؝��/'�=e�vD�܉(��I��a8Vo�y'�����nb��xCu/Vr͏S!ɹJO<����w�P����JJ ���j;|3���Ⱥ+OB�j�ہt��1-���c�R��q��[j>��`Ө�4�t�6<ǥ�+��KUއ�s��0T23�3!g��O{�)�"�j^�B�e[f���U�S|T)�Հ���A��H��<MHV�V�:��@�Dm�lIIW��x��)g�@����?�
鍺�Aq��RC�-�;��u�M��w�|Gy��;��h}��gd��gJ�a��R0Y��B2�������U��7������Xqf�P	5��DhY�0�ʲ��l�'	<x/xoe3���jos�P�e6�;��e��|��m�����2�<�U}��B�$J���')p_�� azP'�d;"m�z�����1����ԙ�H��7�Z���frW'F2vͦ��2��8������Vi��YÉ�v�5� }S\�Vc]����v��&��K"��0[�=�A:��3Y)�[}�*�q�#��Ѕ��+�$���d.����;JQ���!�3��g�%��~�X0� ��]�^�$pbؿ�'�I���/��-��p�� ��q��)�7��=�1�b�Y_��q�`��B�1���ٓ2Կ(�����''�X%5�|y}vR<���l[��9����}��zgH;(���� *�RT��� �kz6���3)V����"pI���n3�:��yga@Wt�d�}�fY�����>�Z�-����w2r�uV��S)6yB(Bq��� �]�Ӄve;,#-����>z�3E�a���� ��*�4F�����@ɶ�u�}%����"&�����EB�0�"dMO��*�P]�۝S�%4��S�O�����[��_x5��lU�.���Q�T�;JS�0o��E��F���2�Ǘ1غ�*�L�$�����f���s|U�WGy&�����J���Ӿ������ZI�s\[Ͼ���1c�b�������p[q�)��,��'�t'�+g4��?lrF�*�3�:``�<Sۮ��M������C&q���K%����)/D\O�i�e6��5��ګ%J�!V�YnI� ��,z����D�}�)�@H��-��\�H�P\�(���+�<d��^I%|PR-����|g��j�3�^A�`0ǘ��w���>H�x��,�O�8R��Ź���Q�(Fu2S6x�Ք��UG_��Н�7c�����G?K�L �뒤�z�K�I���g��J����Vʫ����vT[\@] c���O^;�c�Fuu#8t�*Ԑ.�2�畎p5�n�߃�������G+'`_g`���l�( �X�8�zG�:{����{���SE�R�¨��%ԄO�y�v�_+�.I
�p���jHz��2��D�)l��L�V&�1I�vMme��ħ�\F�E�k{�[LkYU^3uգ�ۃ�Jt��靮������NH u�0,�H܉0�e$�J���$���i�w�����A����9Bo��n҃����0GD�}6[�gщ��e��D~�TKZ��=WOX]Z�Y+�bd�vJ�Ng�hٛ*	n�(͘��#� 5FP���!0���Q\��"��y��r�;8�`�pN< \�xM&�	`�e)�������J�NA�V�y����@	r8;�^oZ'J>F�R��x@��|}dN)�.��u�ބ;[�W�\p��裉Ipho�:��Wۙa�Bkǘ\�G�`\G�#���&��o�$�u���Q��D���5�UP4���md�:�(�94�*<�ֆ{Dm�}"���8����փ���3��(�y<�
22�yZb;���іQ���{j��`��u� �V��r@Yp���x��o_ENa4�96�IC!������'�+�ɋ���ʝ�#R&��@V����V�-�Gc���?ɩ�!ǫ�Q��B�G "�N1��%�&zY��D����@����$���fTfá�-ei���(�:�K*UY�i�����C@ਞ�"+B���>,�f����m�3o�$�w�j�P[MkB&lj���`7���x �Aʈ��xK�T޶��SG��������~Rж�KB�A�~�L@�����-�Sl������ ��"P�Y|���\�o��ooł��.��O6Sm�w�S��Y&x�GId��'A�Yy1S�$�M����a�`���Zz�,m2g�i.���f~��='C[.�7_c�R�q��c)I����$��{@3դ��M���l���L��Pq�X2NIK��T۹	�W��J���������)XY!��Q� 7�vm��%gl1����rC��_��Q��0�k�b�?�E{*�;�n@��.��/Z�CC�5oX֡�d��qy;��&iܠ�����>M�.ƪ��~l.�L�v�p�B�B�.+d�J�U���e�,�X��B3�P�Y��2�N0D"�b�������0M�o lϸ+���V,=����z�^�����P"Л��U�TȰݮ�Ë������8�����I2[�p���D�3P,�@�kt5����6�PN��9ː�7A�b&�һ��`M��	���Ղ�j���3B�O���D����.�( ��C�;$�DD���K����x�đ�e�@Z#�/:�VA)��D�*$�����8C�D��Z%�_XuU�c�i?(ir�y4|ۡ��Ś��@���(�-����bH�;DW��t�JA�i��j#	�y�tZ�'֍~���+�v-�e����[�-A3���X��H�Np
p �dW�V�'=H���I��8f�a�h)^�>.� ��;`�sA�t���)��X�+6ϦS��٣�Xu��Q�n�,��ہ���"yw�@��M��	3�jJ�܏Rg�sLөV׻���:���gm��Զ �� �-�7}G�V�Yڱ��ъa��	��=xN��r�?���TD���v�:����s�WEp�; &���QӓD�̱zg�T�.H>Q��E������a��	rrG{D��C�������x'��m��������7X*Ɗ�`Q��e���"k��-?��������cB7�f�/k���M�M�K�q��ʲ�>�⍃EEt����T����F_�<�w jcQW���Cq�LC)�b\H�{ ;�h�"�f����|zrG`Pش�����Y�bTҲ(��@���$����a% cZ7j�7\Aѡ7	�5��2��_�-�����E�o�V@s������HTu*���EB!ߠ]g�X�����;���_αz��s�0���_d�A��*D��i�BI=F.R�"��g��RQ,w���
9u��`2�����P�K`�A	�Z�$D�"^NV\g7�eq.t�~=G��G@"�8c)4\�-~�ܞ��kN��p�����0�@8N������`A6�,�dO��<�A+��	=*����mm��T3xR6Z��-c�1�����yg#:7B�44��w>��@�ڋ��X9@~��4z����<��|#�ӆ<M�*�-O��?�r%<�jO�d�תJFȗ��s���:�1&� YC�ܔ��^�����YC��6�U*�S:Jp���(b�ɼ�����r��}�U��_+�oY����]�I�"�e�y¦�!Q|�+��e��X���މ-Qk�˳�X	dT�]0�����'��	%J���\�B����\5cȷPŒ3���:�V�5N����dM0���W�ib9"�
��k��EE��XusI4M���z�����r��J�s���e���������݉����t��r�	�q��$�
m�f�x-�E�]��q�u̈́��u�@��&�WG�ͅ3��V� ��$�Ƹ�ٿ��)���-k|�j�JA�11��������8�c��'�$�8A�S�gϳM	8CR����|���k�òi�$��+cqe<3��o]w�+A�B�{%��e}a��-��L�߅(��ҕR.�y��S����v͟�N���ka�*N�u���<�b#�ؒ4L�̑��X���fR%���
�$'K���u���/%��O�9Uz8���"�]�.��cz�$��Ш�[wEۦ�!r�ض��߫aJ�Պ��u`�5�g�oR$���� 6ᶴ(b�N���ߜrt/	/���O����Y��s�cU��g��ճ�������k��(�K.�p�!0����/4b�W���ߍ�R�ȇ��[%�
�[K��*�lē�5���%c�*+���G��}����/�<3擉`����#�tS�9����u�f.�`�F�"�(���i������AHg"�2�|c�/��Qo��Aa��2��1��v4�Kz��xZ0�����U*+��[�۱őXR�A��c�=�S`e1����x�F-�*wX�Qg��a�еPf��{��(!|��n���M�O��u95#�ޢ��#I����$�aE2��'��Yʩ�c���P>��):�[5�� AI���1���	Yd��x�$-��_/��y��y}�XJ�^�nz�ϥ$��&|�_L|Y���e����[����Ob��A���>�]O��Ж�L1۵����iK����Q>���5lG=Lv9��e��MW�߹I��b�`�Hw3@�?~��c2FȔ�{nBV�%���/m��ㅌ���Q3}飇�טnr��A���],��C(^��Wyut�q�i_öN=�ys~"{퉀�g�xs@n�.�򆭮��CM��TT�@Y���NZ6��(z(1U�.��Ϛ���y�����Y�b�v�3���uԋ4B�͌y�鍘�s�^3W��4���I��S�2Y�h�X�0++!�\\L��֛C�����c2e�B�*jԪ�glC���Xe��j�ZV)�����ٳ�$P,�e����s��1;9�m���B�]
3��W����En�����%t$�}�~J@����%�����gJo�]��ۋ�;G�p��}o��Jk��F���f!��������u�N2V��%=5rH��gdī߇
6n���A���X��H��	H#ԓ򽠖]����L.T%טF��_mF*����˰���)#?I�U����"�E��zN"d|pZfY?��户^���.�������ͭ���z�$|�#�MvRY�7KlT6 T��@)&�st���pN3:��^�����6ܚ���g�����ĉ�Gf�qk�Y� �$P Ҳ+���&�oC)��q���Ɔ�#|~�j��r#��q7����?V���|��>nyh���H^VXnII\����@���!|����(�e�]��|�Sė���+�+8|��G���U�\���T)��{�����+�J֎g�A��ϡt�C̻��z偨Yi4��tiRV�Ӹ��g�)�W�pI�"l(k;�6l�pF3+�s��&�ե$,7�k�c5���u`��PlSD.�W��"يr�,�٪��_��YQ��փ�B�P�*���I4b�ӳ�nlAqz��Sn��z�C8�<rq�J���`��~H��N�B���*pm˕
�%MLf]��?��p�Ձ���L6�Yˑ_���^��$־�́��ArB�'c�Xiq���rA짭�����B�� ���C�~�`�;���a�-��e]f����%C��]�|D0�����\"�D=Sg!�p����Bi4���J�����H�P1m��������̗?M��u�*Ho���91t�\�����9�M[	"�6.������5=z)��y��Ӈ���0�uq��@4pA�f.U.����$����k��O$�wݥ:�3��{X��4vX��Zl}�n��#��$���7v�"��/e��z�os��l�cL��a�:�Z�y�9N�L#�;����P��3�eXԮ?tY���IK�n+�i�W!�$�A΁�u��c:r%~�_��E�ay����qN���C_q��l2��w��D����]�sڋ�-;�]�yVF�K�6'�o�
J$N'���ge�nj���=I<�ͯ�Ai�v~R0�L+}>�,�x�쫛 5wH����9�Ua"�F�d3���W�o�JZd��(>�@ ��ٓk�ѥxZ����E:Q��動kU�_h!1l���_�Z�B���(!bq���=gc�ʀ���?�H���2�P�~۽���i�uk9Ƥ6�"�L��g��߶���AyO��(,X�?!Pp�	��b�9�4��D�yH�s�sғ������Lw]��p�)�:p�4�q�A�53y������hDػI�n�lGH�g!�S�K����9�l�5�0h|\��Ɋ*(*=��Q5����sYL���џ.[��`[����󛬅~����H��}U
�����M������"XB�A�{�C��X6��u)��X��+:H�/PMѠ�!Rd.���8q4��JQ�0�����Dbc�OA93��LFq���Ō�6��R�9���;�����%��He;z�2�t�)BF���蓡���"B�eU����ʌOBi ����/ar@H��DVDkQ���UX�T�N��P��0Z7�5@�l�H�6+T��?EҞFnK�ܹӑT��'���& �*��,M}σY��ARu��A.�t4R��w`�;`o/5ƜK}zGI�r�� �*��b�v�86e�6�HQ^	L�ʫ�pL���d��"!e��R��u��oW�i��g{�1B"��� ڜ��J.2���'[�3Q�#�ë�.�P)"`5��0�	D0�` 6<�:i���5]^��y.[=G{����]�kx�@q`�1`b���.�TƊ�A�r+6���`�n� ɭ�8���܀:�D6̞�k6sB{6w�!\��1
�3���7S�yq���������dَAL�Q&��mlޠ2ن���#��P���R)%ù�&�)Iٳ
�m����!Mhި���g4xm��v���?RWau��Yhk�x*�.K[BՏS��ǓX��kmW^ѭ���������!�AOӗ��#p�	S��z����jU���[�mL Ⱥ��x�K����4�򤶪fp���c�Z��| ��J�����9(��7.���vU�Ɇk���M��<�|5W����h ��(.�e��\O�/e��o���N��&���i��D���h�cq4�1V��ɢ[�`Fwz��;���_.qc_�ؐ|t7C��a�Ǯ�䂎�{[;��lҫ��x:�R�ҹt��q���"Js�k8u�M�K��a�o�۫gq��%�w���Jї�_�����\�>��n�8�iB
�1��#vE�k��^u0`~ޒ���hG1de%�;�.�N]B�s���m��I��ŢC��]G(����Z+�^�St*������4��[����5�Eh�l�J�?_�#�iUx�=aF�^�Y�FZh�	!)|l/];�(��b�w\,U�e����"�na��:�+���g�KE��ЊG@��DA��'���H��IdE���K�����r�͉�{_G�BSZF�`��H�KyFpZ�䖃����\��d4^0-�#��a�+S��UB��Hk7��\�w,q��"_��+�n��)��.�S�j��Ԭ)�����sܾ+?��q!��;`%{�
�0�=4gB��*D�Y�C����<�N{
�y��*+��?���C���P�P[��?���O�n�Q�`�=�]��e��$��?�p���*�O%�W/���T�+.i.O;��.J�΅oG#k^@��/�K����QubY��$�U��P�ٴ�O�\*Ȓ�5Z���"�0�5/�(���Z�{e������O�5�����<{��HjZ�wO��E���V}q
�i����rU�7j3��w%��8
P���(�/,q����ھ�@?2��V���J,:�_\%�Qn_�bM��I0�
�]E��Ó���B����;yG����6O�%,��`/�^~3����p��+ePu1�h��[>7U�;b=y+���v&�Qݶ
�r��Nd�ú�C�h�r�68�HO�C����AaKt�Q�5�1�s���E�V����� iچ���#�rf�]��b��x����E������wC	�w��b����@�X˽E��<j�xuY����mq���r�@��T�@t�_L�+9��p,��
��c�6v!�-ɼ�`#�]U����lI�l��=4�X��v*�W��LNؗ� �����\7&:�t�ɂ�B*��3i7�
G��)��j�9ⲵ�b~Μ�L~��7��^���P`m��8���NÚ�8��	Wqq��×4���==(���tC;W�؈���U3Xy�=��Q{5�����gٌy�L���0��/h��6�*��9a��+���ԕw�Y\螵��-���l>z�t���o�b87��'WRy�P%Yh�5_
7 m�P]4QyR�BTEE�Gx�ݓ
� �;%��W�Y'�Ϛ'H߄�jòʗl���$Ȕ�Bw����=T�M�җT��$ta���^�㝾��
p�C>g�{SH.6�����<���{���m�φX�&q��^u����*�va��Ē���Ձ`���ܶ�X)lpk��Ce��B��l���n�R4�L�⤈yԵ�G)��hhW��m	G{�:^��g�~"�a�
>��ˋ�šs��d�C��D=�?���#!��V�?S�PM0����%�,=��-IX���.�t
]���"�Ղm�h�ú���[&f�0X�������*J�h���������Y�w��u�O�{�t�[�*2"谽��q�җ��:n3��l������q���?g�܇R)���j��ڕ{��0a=tW%����[��f��qI^���|r�ɲ���`����Qy7�P/\��Y�^�׽"Y���ˈ�z
���J�����8��*����<��9F\�=�!�G�����f�-��q�0�f�\�Rw�A�0�u�]`�} h��ތK[��&C�O�2?İ�l��9c��������Q�:�D�5�?���h�UDS��畐�,�ѥ�\/zB-�����Q��$��뫄s��N��M[�7���
���"�P��5P���Vp�uœ�6�uacٞþ���mB)��D������9�i,���*L5�=D�K�f]#�C�?�����~(0�c�$C�V�і��f�d��E��B�Ge�L�������}�g�Mᘢ�op>xo9��RN����MN�.]fn�f�U,��_�K��d��B�r8d׮�,�p����۔���;1���I�G�Q�ĭ[�m�UB��@�r{�U���ʶ�aO�"#D�G1��h!��kә�D�A�g�~��4�՝���G?3�_{H���{->?P�$�?5!/�R>x��l�!�<�Q�� &��Dz����^x��4#���3����.p &�PNǀ�B6	��L�C�M���2��ꈇ_�9u�Hm��ͱG��A!Ú�M��������12��ϖ+!�-B�✻�2�t������P6�Y�I�Y�\�^�X��+;u�ʆ��t��`��.�M�?&M�7ȿ:�4���eӅ 1�������mǰc1���d�&��Ã�fl,U��kRI+,p=Tr�;�W����A��!��	��3;#`E��
ٰ'�7X���Ĩ�"�HV��
J�|Q�i��m�r���*Pf�L��7����/������H�ŚH@ԥ���:��a�?��o�Vvd�\pXS.N�1�L��[���e�� ��o�,ݥ/��
�cq������vCMR��An����ޫ �כ_�#Hb����C���T��^7����2\ S�9Բ�=���$
:
�0|��(&� a��W�e�bz'zI30H�\@�N�blQ��\�^�����)�{��BT$�m��Σ	�-��-D�R�	�fĿ����Fwص�"tsa�=�Fd�o7�5����P�X���H����/_�qw�d�����t�m=y���rO5�_�1�(ꚶ���8�i��X��s3�����40E����w������J�Q�m 8�L��$�?��Ie�\GY�F��M6D�	��3\��*��*��$o�>�$Q � (g���à��Np���fQ�Z'��OU |�ty�ܫ�^[`c3��/-��{?�s;8h�����l�e`����㪩�?��1����tO��v¯=��U{�8�����3�F5^I���q�$�ͼ�%�9Mԃ6v�T<�E��q��9�B��%ѵ�u� 3��� ��O4��bh�p��Fo6~2W*f�I�4a���+��Y_i`��[$�+�H�}�� l���X	�>�]��M#u�/� �0�_紝�.o^t����N�Z����!F����8 ��|�]��t;��kZ�j�9��!��6Dɓ[�ݸ�'�a/��Z�u��(�k^��\H�P�<!"E0Ը��)���Ax�6g��ew�3M�wn�#�m����%瞈�e[ �ѓL�'yN`�#��d�8L�ጜ�	�}�yN�N�#��B&��əm����ŉ�Mύ�eǂ=@�M���<�2��t#н���6������@��!X�l����Ӣ�ֆ%�<�=T�.-�A�ߏ�{�6��4��*����G#�ꕸ�-��1.8��Rhno�J������̺$v�kI�/�?����uz�Q�9/����E&�J.��Џ1����N8������R�hfrNJ�,�[��,�E]�(�EhX�.���y�� �O��-��`�:Rl�r{�{�	>X����'����4����#v��\����ao�-�M|��b�AD�h���ۀ�ߜ�T����P�C����#�2~�ڕM'xY�9ǳt��YQ����K`�U�zT��+����,C
�?W��>� 5B���T�	���b�;2�ѧgd�z'��Ha\ըƑ��S���h+�Gi�z/;ڏv-u2����w�y���x�%�-���/��Z���.WP=R� ���k��Ck�
gt�u˒��JW|Z}6�t¹eӺl��'Г���GOk��q q�,�����&\/l\���\��ҍh�,�o��I�����
�Ϧ��lz
$w����z�֜���Zw�X9K��7W��l�0&!I�)���8����O��x��t��d��h:�C.��!�$�9�8�9Ě3>ERk��֘V�*q������p���1����Y��A�Im 﫲F�����:��2�XV��R�\�g�5��~��ey;��c�K丯n�2�3E31X�x��X3�I�HA����8��\)|� ����o��d�5�-��H�M���bW���PA��~�N�KG3�#������dٺ�$��R��&Z�����pMj[�����������,7��<��~zO�������ɵk���V�����X�?�3J��V��9O��8��m?pkL�H,���nXq,(hc���s�O���6��� 4��B�4�.'����U �,4U#�T�����4	�3�5����!o�G�;�pTh�XI�3��pF��ڟ��a��C�/4C�"�*�/���+M(��:��C����X�g��� 1-0;6����;�\�\wj��b7���kD1l�4N��� ��#G��إ��O��������	�;bƍ�N-z5�sDYPӇ��y��.�nZ�
I�%��;n+
[H2������Q�((~��[,7�~���*�\�"�΅p���u(9Q�|��� D*������*��㽲^@G)�`n�^��s�5J�%±&5{%h�w�HQ�o����;�����׍9�X�b��&��	^D�1�j4pa�2�7�C#U6�H۲���7�l�[�_�0�n��"Ц'�c2��j� ��2��z���;&?C6�j��h���}�"v��<1�R���~���<����H�nW�8��ѡ�xt\ڎ&.m/6f�T�\1����6�������M��d�M���Y2}����U߂4���$�]yp�ҴՌ>��-o�Cn�1[�y��4����Gm�Ŏ�N|p�_�T�:���~Tb�WU�@	��hU�6�Ҳ�?[�$:�Nm	�_NpC�^�����)kjc�����m.K��Ǐ	g*�o,�c�0i���NU	C|UJ�d������ȭ���F�g>3�k�8Q�{nѺ���3\U�4�*51�Ng�p�^��4�֧|���(Lf�-#cM�яLU�w&N�e�vlb$�a�Y�ͥ��7�q��n6.�G�G�=�*������	�+����^����p>��/�=��N��P�9��Ms��Ѝ_�����MG�÷��O�~8�v!{�.�`{F4��	d��#���.���	��F����?x8Y�2�/S�2��_����#y#U@ ��n�����H�=�ɎtY21�	�����k�ｭ�dy�6�Z��
��G$t��<�"V��^����3�K�_��G�&�n[�K-�#̔���.��!\�R�U'��y��}u!�r5���`��f&)E+���T������Y_L$����N]�F`���iK������c ݤ�L&үV8�r%�z�mK^�WO��q�T� �CO7�	h����N��p2���tpx^��$b ��7��4��N*o����OI�������F<�w���t{4O"���d�SC�N��~��B������np%ug��Y}��SFN�N#r
�hD58HPu�I��#�@zsH�����JŤO�2�9�_ ��5$������ɧ>�i�Pֿݢ�ǋ�tP�H�<k�25E>l�TJ�
x\���l��.,b���<��Ȇ��\�E(m �^R-�	FV��^��YgA�Ŝ:'z^�ҭ������d�/V2FN�$ץ#��{4��� 4H٢+_?�K�hL����qp^�����-뚃�+��lr68�K+ӌ���
&���4�;%ZN��3��3X|��8��g�*���)jC��$�	qe�
�a&����,Ǝz�s5!Ao�G�)��s�Z\�O�A2_�W��l�H�:F&�(ҝY8q�j�I�BB�,���
~����K�><��8I���%��<�0c�N���d�h��O���Dō��K�a�>�(�C�S�j@�w�%&	�����3B� :-�a� �U^����;tX���PS�s�h�n�l��<&�yFW�n���s���L*dP�7Z���M�E�w�~�T�Ҩ]\���.�)���.���-I��Ҁ6k8~D��bw-8ߤ���� ݂֤�9�ݿ�����@-(g���6�+��VێIg3P��>`������k���z����/�����]Hip�r�[3��n_Tzl�̧	�&�R<U��ʟ4&�������$ք�{x5���� p��A�>xZyY�c�7<��/$(���Ј�F:,���#�,���F	Cqߑ�OoA�~��x9�lt�]҅C�|��IUr��bB�3�ǅ�7}`P� ��}�����w��a���Zu�ԀaQJ~u �ӊ���w\�#� �J�"&��]������֠�Y;�\�؂��p-����M���]�lZ��i�;D�q`z۸�Ѷe�J�ˊbm9��_D�s#/x����U����9G��\	D|��L���Q�-�_&�?��@*i�s^ʽe��,:?�n�+q�(�(��8�j1��	���*�&׌���=�Mʧ���`fs�K&,{`�m��{�/>��u��h�6�rz0͌I���M\�-f,���Q�&�vG�|s����V�R���Q�e����3��)��v�~\�����K�qΪ7�k��W)��Ql+�@ʥϪ��� 7_:J
XɢuL4��^���R]Zw��+N���9Z�+i�܆HǕ�oE�*茨�*w�-�0�\"����J�J/@)��̚�����9�������g+��!�.!+����8ޝ��ʡ��١��N0� �vr:�,_s����6�U�)|�7�G����QP�ֶ�*��\_�j���36Q�8��JVZ��IGq���b�q�]��DD�*ü�iň#�������ެ��X}|Ih�e&cj�F�e@B[��[�6��Jif���#����H����x����9~��
����N)t��Kd.&5Qn8�.�ۈbHw^�YL���g�(qݙs��s�$�?���rD�/bY���zZ���j���6\G}+�N�07,���'�}�K�eL��2�?K�Z�\b�� 3�{Q`G�����ՠ�mp� ������,��뺀W_%�)�$^��ݼ���R���kyn�]E�bfi�?�����v�����
�ґҸ]�ֿ[[!e\nk5����%� 4���r ��`ڙ&����H�\�³�3_u�"�?l���I��#�,��ȵn2�@~���ԋ7��\Y$h8��R�I������t�x�;k���OZ���]�,۵a����K��_T����$�������"�h�1�sن0���{�b��̓�c��n�c� j�.�8T��s_�t���.1��n�H�����U��.�̏V;�����%���%�TgbVY�����o������o!�:�3[1-p�>���[���{�`�	�*�x�s�Yv�p�o���.:��?���_2�p�p;�`\�\���Z�� oF/&x���Y�Я_V����E�MQ[?Q�v�g��KA'��W:��b�Y��=���x�����E�*J[�g��`� 7��-�I�N��y�3�%'�8O����~��vƒ~�?�����OZ���ɇ��+�g�}�.<�0�
��O⯭��i�C}�%���J��G63μco��=���W6�V|�J�l��T	z���X(o��?Du�{�?{���K�m~�� ���s2��-1lW�\�18�+й�*;T�M���[N��&݇�?P�ֲ.���l�0|���c�?k����M��;�Tw��!��c>�\��?� A��Qeo�GGZ,^'
R-�=��SU�v�R�e���*��OMk3Y����96K>���m������7�u.ݢcx�ҥ�+(�]���L�Gu��EA�"�a�O�D�r'�=!�L,?��g��+.9"�fﬆ^ˣ40:�7�����`�B��U��0�}~�ã��v$R����n<1UI��1Cf�q�
S�!l��L���m��/��b��\do]קlϧ$f�6
1S>WO���=�pP���E�O_`d�s"�Œ��+�}������p�U$�)=��|���~K��s)�KNW���h�9Mv��zM��[w7Q��I��fY�o3�����L��\)dX�!r�n:%� �[O����>��̯'rh���/s��C��)f� N��'�C�|b�fwp؝~ǕǸ33��*�YUЀ4�0q{A��ݍ�t��𞹾���"�������餡u�۝�xg��s��nP�Bɣ�����g5�lr����r�}֎���bŕ*�Q)��^�NoX�m�q�.$j�n�X_�Af�k�y�Yt�؞�uVBe6��L8q	�!�� EV�A�,#
���`r���Qɯ�N� J�	�{
F�;���ٖ����ۯ��n0O��<ׇ1ü���R�SPfs<l����l�N	�^��(�P�� �$Q�ݘ�e	
���,�L0�6����I�J��$�Aɏ��/�-I�f�MF��9sf��$��N2~�"�
䲏��9P�?m�a�8I/�&�9w���~�Yhӭ5�(���	�pF5�p�F3A�N�1s]q+�-�3�Փ����7ȈK���H/A��Xe�,�z������?�О.�
/C�*���@�I)Vj2�O6l��$��������N�i%�y@i�-c��:���K<��̜j�^Ŷ;��鲜o-J�X�#�/���rh���[("�9��{T�b���Xo������@bL��[����~Ե��oŝ���ǔ7� 8R*�5�|��Z�{s{9�q�Դ◴��9Zؤb|���RPpֺ�<�\�ɸ�G�Яח��_������֜ӳZf��R1~?�x��"&� h���!6d���*<}K����\�2Ob[A����6�,�g<l!0����:ꓣ��{�X�V��:q%Ł&ti]�Jm�4	S�:w�^��>g����D�fr�n�6	���̉bqc���i�FŪ�n	��g1Lo�ߚ.xq�͇s*��=��7���5M��S"�|R����� x��Y�g[`���Q�.���[rs�8I�=�;���&l{C��k=�󶹠�s�	�K���=N�'�0`̱W2� ���6��Qhu��M������F���o�P��o?�҈c1�3	�����)�h�����K�����c�W��4NΞ�'��j��� OuKCJ~�#�,^���I�� �PB�r�dT��ѩ@E����������mʪ���O�%
>0��P����%�B:�X��B��U��r!@;^/=*� 3���zڲ3�[�\���Q�X�sĲy��	K+|��B�2�;�� �*v��:/}��
��cc��g���UKc�brͯ��^Ŭ[h�:a��Kuw�2�`�U�xv��+���C6#��T.�l��]�j���Qk��.���2hg�QJ΅�]�[@\� ��Q�Жۑܦ�L����Q8j`B��'����<���l����6�rJZ8�mb�F�G������*�W�;��?D���