��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�Oo�X�=e��F�O����
��X����j�ۤ�POd�x�t��?�b�v�JZg���d�o� g���x��ki�g���h/цƴ��g$�Zjg�=�?�����J������9
7��%�r�N�q�w���zK��� Є�f�l��(����I����}��n�?�.�w��o#�k�c�����18~�_�w��L �J�Ae���U/
�|x`q��[ӁX�Q&Rc���e��)�W�M(濯Ie���$r��vl�����Ɵ�1�`]l5�3�Z?]�P,��V��T�D�x;�(��vf4��=�>9��Utχ�h:��I�m�NH���k��)���T��0���G�GG���V�	b&k��n��_ml�`����b"�s���Z�����2����J�[�n$�[�Y�R�w-iILe���)q(I�Gr��o`5]~��F�uF�l �"�����~��.��JzF����#�j�H��z.4��h�X�ē_"(�&�XnA�w�h���l9Ra�u����_�Pzl����=a>w�A�+'k�f�~�;�،O&�ړP��"�j��G��(�3S���A �[ĳ==Ŧ��-#k�K�e�IQ�|�݄70�{2O��Es)�@�b~3Y�v�q��Vl���:���#h�#}����ia5����xC���^q�Lk�a8]��+H`_N��et��^�C�\1F@�@��F}�5脓�ڸf1 �Z�� p�E��Jo���#����'�7��D�z!�T��q@�$~B�k\����W�m�]Xb�B��vf
b��}5�; [�(�sS߽��ɂuv�諛��"����iL�������|�tB��$ѿɾ2\)�����m�.I���#$ �:�\�Ƀ}[�����o鎱�M�K��}�#��rE������*�V���hO�~�й�n��a�Ψi?h�pt�m�V��f��Yz��@Ѝ�̈́�9�4#_b=w	:.���-�ɶ�!�q�Qb���p�+�ӏT�������9;3I"�a]":�*�xc'9g�S�t�h�?��?��IN6�G#u���,�ʣ�n)B�.:@���sZ�M��������DS�(p�zi�!*2N-�o86K	���c���EG���*�d��lA��o�H�s�|NL����2�q��Fl�6��}��0|�W,l"�%j�V�l]�Bx���1�b5�i�������|�-U�ʾ��������:G"�990e���i�s(6��W�)w�.ދ��F�p����Q�*�<Rz�Y�G[=��7�h�����7���3W ����_U�����R��=�1��u_h^)3��� �(WUѾ���oP+���U��U6	��~+̻��
`<�d^@�,䇶�����8ʍ\�M-��� ǟ`V8�P[� И�B����aW�}[��]�)��Ӡ�h�輷����6Y��1�G������
���r�0⼆��������٘���sb�~����U��!Oz�]{<HG�G�
���5p<�!�zf�C�)@0���8d2�(�X�֠��@�u%�#ZM�8S�ޫ�'��m/l�	s�J��)a���ӫ5S0w���|�#Hs5#�����S۾�;o����"9�Y�T!R�M-eQ��h��0 .d�'�2Fւ;3��{���gÃA=��z�p�0���q/�d�Z� 
�z����%ó�q����y�?#-up9�i� �H̢6E.�Imi��K.�-[N��^GcW�a�����l����^��9���us��߰k�[8"����]Ǔ��Jj����$h��ߏ�ͨ)�m��-�c<0S�M�/p��b*��Rf�rzk��p�H�(D	"��d1�gA��~���*Ǥ��C�=O޸��F�Lx�GBI�M��wS��Y��&�*���:5����P���E��vNd¹U�mh���Ǚ����_:�Z�R�Ͽ)���7�Gw�k��{���U�;�Cȯ�6o;E���~���p�o5�aL>�f�Z$i�jn�vJ�$�J|_bh��t��N���\� �	�7�bE�qPN�Ʋ�:���JX�ķ����+.�[���Zq��P��1��U�G�g(�}gF͒�ʴ!�Zm]n��K5b��C�Ҷa�d�Ҡ|�4d����?�Ò���L��ܴ��G�|/���5��	�r*K|�M޼���aj�\���ڸ)�ENpW-�_:-P�'W����Fώ/-F��zZ��?��/� ��L0eALQ����oJ���[U{|�񒶬Tm& �H���GU��5U-?��5e��į��0�(ف��K�R�z��U]�!J���B�o7��K�
흿S�>ë@d�����P���3�je��'�I�'83��K�9�W��ŅӰ
�t'8��oq��uX$-��)Uv�Z�|o���lQ���39ԥ�4�|EI�IAB��a���r����vb���wIsDr���ƣiH�Ҷm&���L�P�B���vxK�	Q<�Q_D�F�*�����s(��g�s�(H�~@��qꌌ�c�Ge�$�ҟ|��ek]r�H&�4FG���&b
�~���ӥW>�L�
jV�uޮ~7�$��T�$�$��s��>�c{Z�Y�8�#7��D�ו��t0)�M���;����7
���	pksk����������g{r~��2A��'*��"��w�m�ݺ����e����	�Ng+�E��ꁬ�G�5�Q��ղ�L�Jx7���b��a\7�E�����an�k���d�]n# �f�-(t�o�.A��5=R�=6@���ň2��p�C��V�B&��E�0�	H�� |�FρU_��5U,y�,��^�ާ�yhh_
S��j˼�ĲLZ#7� �C�C^~v�6���M��:�X&��:#�N��ş������������m��G�|6����~S2#|�'�KI��.���|�������4�~Q����yF�uk�{Cdp�ISY�����F:E��������RC��ou�k,�m�n2j����h��2-Z�2�@}kw*I�-�J�s(��ε��\��£������B��(XJ˞ϩ$aEtN���f�K$���^Ƌ�qx�;z^G�i��b���7�ԯ�@Xё���l��u!�s�LU�x�����i��"<�|O��$��@b����f�Q.��F�R']9��iJ�Y�m��v�xdk���g4q�Y�Ų����\ZwPw�.�J�[W:��;S���4J�1f��v,�˰��y#����*� 7�$�X��m�A����g�~�]ߤ&n��r��)%���R���A���-��)��	v�Շ�/}����t#'$$~~'�u!�K\�I��_A�Jv��k�BRC���������%��Q��*�;�C���^���!�+��(�@>#�>�HX�%��_Y��(Ӯ� �Z�~�5]E	;N�%��~�CØ�07���lSV�
L��;Y�����!���C�X]�߉2:��G�}��G%���s_�	�_
��j>CG�,�@���,ۤH
��q���b�ۊ3	kk�/*e�AT�	�M��`y�Fyݤ���P"�a��`�6d�[��Xq��X��fL�����V�&>|�8�{��X��d�s��Ʌ�Oy��!��=ˁzD�c�0��f���sB%���/JK��y/-���w�2���������9"j1��f��Kp5��Ӈ�T�[�	Ei�|Z�gvwc�}�&~>���l�$.�٠%�Գ[����4v��O�}����O�̪��ɖ $�w�'��68�\��H��kK�(�ʏ�~�q�|�9�/<u=�%�ҷ),K��;kC��<��UOi�:P��WF�0�[W��e�������s]�oT�W�Y�˻@��-�¯�C��va�N�p ZP�7Is��:�%`� �4�v]�EN�1�D49�5x�$��
��;u8(�rA������এ�+���y7/w��b���&h�.�;�5���I��O	:��h�����]����n���	���ȅe*�����(�|P��׿�z ڍ,Sy(��Ɛ��R���$�OB㘒�C���� ��.��D�x��0��#^j���>����{�'�oT�T���b
*�0�R�z��U�d�B;$�d�0�����/�f�Xx��t5[$7�g�c��o~^�ij'���|KY�K;����O]����������a�v�K�|ۯ��C�}��T��Ra�V��m������7	q����:�吸��G�+��UƓ~t4��!���c���)w*��ms~\IIo���L�&�:���>�Vg�!gEn���Y;�b���/�u�@�:i��ⲟz����L�ݚ��*f��� �4�������.�L��9��܇�).5Ɏ9ē���n�*i�>f��g�Q*�]�%�����'��φ�:���3��j�Y*���f��}���\/����Q�b����;C�S��U�h���V�4/���Q�^$�K	������h�>;B=y�U��Nw��l��J5mdǣ������������PX$�8�Kw�GQi�ԏ:���B<����T��?9��s��8�`�:���_�$K�%�_�>�4Q���� ����xV���Bꕭ
O�fJR��ה�Tí ��j>-Sѡ�/�F�)|�f��4�������Tf�������t�����o��066t��ܦ�.O��m'��p�g�ʢ0�����*�8P��<�O�rא'[����0u�b�v�:B��Y����M��2rژR�J��t�����$��R���V79C�oH�Q��R�\���N�) R� �d��Bj�5�xϼ�T]���E�T�mh.H*$V�lg�#]��LTZ�ǟx��bU.�r�Z}�l���BK�4���I��>Pb�O�z2^h������"O6�w�=�DĶ$��S> ��f��=�?�2�����}KZ_��C.������Z�I5��TW
��#zE�vٝeGL�����pdH�������(�Br	Ұg$��3�4�5����kB�[�[iҖ��e4�`����OT�L�[it0����&�<l��>W/��q<и�%�^�n5��mr��� ZNےw��sH)<^�ے��=o�7f����8k���E'x�M�j	1$7za�-��&e��K����$Y���t%/G_���[��q���#����JC�d����˿�!���U���s��\�\���/�Xj��_Z�θJ&`G��y��'�[JOA""�ћ#�����=:�7�ʷ��g�z��M<�p�6#۰�����Ya��V�?wk�"��:�Ꮫ���W������j:������c"�`���w��� 7��%-�
���(�ܵ��i(�4Q��1�{U��\,Ŷ�-|弋�=�&'O��ɇ@M��i�-��g��ؐ��|�>ى��Aۯ}R�=��IQ��9+
��6 1!vJU���J��#09|�.�t�~�� ���M ��*[������T�5.��P�(RՄ#�w���F�-����wL압���ʾ�B8�!ۚ��D��q�œCEK 2����QS�sF��t�8䍰 ���uM��S7
�_�c����7��C^�{M9\Q B&���_�5-x��b8���X� pd�����Ζ��kӉC���Mn;��J�+%9#���
���
G���~��䄩�L���(�
�{�Lx�X�X�����(u�uOxU����X���&#y)���i���q�"Y�6��i��E��cZ=�Q��R�T�"�X.�}��E��0+Ϙ�ِM�Bq�<�����.�H�R1\"� 0;�����U�l���[�C���P��.B����;U���X��9�ŻK��_����k�m�z�m��>w�߿�������|9�#�S��:�1譄z��m�TI|(w@2ʚ\�#-Q��u�k���(*�
��֍W�r�LTҎg=)��g~�<�����K��U_�|%�/�i��8-�$�͇��K��W�+Fb�1�ۇ��j�ZC6��_RI�̖ ���l��
L�����c�J�?'�@-;\�,��&���@W�AWП���0���#[ �[����	_d����)�+�3�ġ}&ղ���Y��&9}� �G��c���O��n(�C�\#5�0�m�Mzv��#Zk4�d��WzNm�H����k�	K�?឴���BI��@�8�����5�v/kud��y�^��1����k��j��K�����[Plqun�g}p�m���zi��_�-��Jf��h���s�*ˁ�J~�4=Lo�	��\��x�W�շ���ic#|�S��֎2s2��ʮ����j��+{ ;�F\،���9�Wt�ݬ�쌦}H�Qz�3ݦH'��DEj�I׶��w^U�~��sO�xw.�P�dBDG���^>�͕M��v�ʎ���Q�7p�}�L(��-��?n�����m���"O;�TTP�hUb����i�OsU]]�HО ��/ι���U���"�>D���w��$��-�%����o�,N�}�Z��އ��g�Np�X�3��nYhLjbk��N21EV���L�4�+!p?<���<)����!��Bs��3΋^�)��o�`-2nVs��Aa�حI��eY�������Ig4kA1v���OQO�gE�h���qɆg�����d�q]�D:���T��x�ԛ�uC���ҁq�vwJ�bVGvB4!��CDT�5y�t_<1���V�� ��c��x�>����2�v�"9
Ckk���z.�\���Ms��d�D�4������
�z����-�8�����yj.B�~�atA�hAޕ�6Рd�2	ͤO�8�
P���~����dֆu=IԑJ��	�z��P�;�S���*{$�y�l�st�"�hp�LdK'Ŗw��5%r�S�����N�D[�*��
�ô]�U�@�F��>�,m�wV��6N�aG�b�� m��)ڍ�8J�e���Gxl�{#�)�9��4Sd72W�C�<�T�AM�Մ4JJ�%��w{J��"�������D[�2wbdּ<�j%����t����W.U���k�z̒n���������P�Os��2�{��/�2(�y-�Z�+M�\T)�J2�M