��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���y�'�>�p#�I���K��xƭ����	4u�ױ�Z�4��  �=w[�5/�)�G��t7�NN
h+��G9w��K��t	;���5k=ǨS/�ֲyb�崜����Hʜxo	YDc1¼A)�YH�e�����T���ɕ٣o�,�v�
�E��.Kf��������s(]��� oI2��Wyv��h���vބ�p�LJw�x�k��Tx���k�׎Y�_�xC����,m��������Dџ^�Y�݂�Ƒo)��9�H����m��S�P�׊�P�
��<_�C|<ދA�t��Y��C{���[���16����$�Iú:)�8M�1���$z�o?����o.W8�+J�0_O鋟$[��k&�z�m��qL��	���u��ng.�[�(᰼F�1����1�lhN��@5m�7���(�%��}�����!b�m���P:�l@�O%4����
��/�Ͻ�i�#�i,x���)�'Ǡ͜c5)Np��"�3�c���'�lg �����-�J^�������	�WŨ.���G�Q�����e�j���nS[Z��u�5)���o��+���K:���BFn��ٱ����B)�~j�*�7=^�������<A�+;�W��	%s�;Ъ���y ��?��m�;�_,�c�vU>�I��*h���MgaO�DK��0��&j��L7���Kϩ;
�]�B%�	�5�f3�N���b���5�ڡ��tN �Զ��$�n�_;���nƤ��j7#F|O���F@N �W��ٓ�>&�Z/���?~��	ƹE�t��o5Ds[�7�"�+b�~-V����V-��"��Ȕ�qM@���6d�gʄ�D�f�9�F35����h�t���$
��'�W��p"�N4����v{V��]�ޯb������ݟ����A&w��48����;\Hc�߫��O`@E(�o����g��߾�	�	8�{s&9�J��W7��2�wKL�+�Mb�jh{�8�"�qů�V��w�P���ꑩz�j!���w�q��*v�	-q[�N겔.$�B��#�M�����
�7��˥'��j�=�o,IO���s<1M�eZ�������X�pl�
Z!�Ձ�O��<@S���K�p6%w%�A�)F��n}��VU�\��r:92�X�*��U_�˩�������w��r�e���Mg����:'I`3S��)��c���R�~ȏ���.;<�,�k��y��̊/�J+tQ�e��V�Eؼ����%}C��϶��9�jPf��������tu�G���c�1���3F�{?�V�(=�E.�]��J4������}�w�&�3���$���h���N���@����4|��5 a4n��
G�����7t��U��8:����ʖ��x����ڤ���G_-�s��Ll�k���V�
�OR_7��b��B{È���T�������G�Qf��,q/�Jf�[GH�F��ZI�<!��90����'�ty�p�G�����?GИ�&xV��W�����僿�<�~��$�$�S�.RYc���Ւi�h8��GX��!*pjb�T9��TI���RؙKlb�usr���t$�Ȍ��
a~�b����r�@87��A�\B�`�t�4�tO�F�j�c����l���3�Ŋ��;zfʀMW�S'�R�I�����D�F.�R�կH/��0���.�]#�ۊ��O���+���[ʯ�I�D��VϏ�ӿ.��2�ZP�r����'�pw�=z�s9?n�0�u`X�bk{����Pm��y%�g"']���7��M������*�7\�v'�ѹ�'�]Qw��c���v:s��!q ��ʄ�ZųH
�3#�uI����X /]��� ��{ǐ�/�i�=�{���4�h??^Խ�[����ѧ��B�6dT��l2.��Vş�˱mqY|��2�U#�n�	'&NF�T�ϋ�1r˗���r�)'����,�1◠��h�H=_��w⻐����S(ɘ��|s������q��)��˅wG�Z��De2�8��;����w�OKI�e��\�X�l��5ӈn�"}�UB�����Nz�0�Y�W%B_L!_�/�DiK�4�	}ƿ�X,����G���_�X��`7F�ٔ�8��
\��>"��&]Ҵ�A���𯬏a�=��[!h4���k6f8RhY���e���ޟ�y��}���"N���~I��)/4�����������g�2h�@���:噽�I2t�(.`�8� D�5>a
�L��Կ=�UyaH��N%Y��W]�ε�~c���{1���~��:)y�z�R��A,�M�%��־Tr���%(���>����`*b��&�lcr�~M�\�y�N�����ߣш>�Yr!�����;%(졼g�/�I�=��#�J�.��F��g����=�	voH��KZr?y<�H�N�_�ݶIc�-�.�޺D�(�^��p�덷�u��� bRE>�A�U�c�Vh9�di�� ��]Wq��ɑ�;��j�D��Fu�#=#��a;��AM��������x�}����������_��b=���f���a ��M��2:�uf�qG���洭�½O�bq`��G*+Y7^
-�ח��4�/VE X'3#h�Ø80�;���}�?jI�C��|��Wo�w��t���c�LZ��vqk$T
�	C?��D�TP��9��ؠE'�|-��$��	<��Q�cЅ|
���.0U��E(�D�/7ξ{�9-�&�[SI*%]�)�����,8�'�eT�q�cJxL�ڴB�lpX��� ���HI���lq�Ⱥץ�����g�1xb�Ġ�ڇ1
� k�]�@1�vC8z`o��I�b��|�`*���|:�t�C�'BȆ]��a�� �,S�5y�6��~�}|��֓]��fAr&�4���:��3Je㥔�/`�7�,w����G�V�Kx�ޟZR�#�Y@p}V�F�Z'K��d�U��=5a��	�P n�^:��w�dY�������L��1Zn���։0A"68��гץ��x��e�RC��y��`�$�"�Ì5M��W�j�-��~�7�f�rgQ�gk�����&5�ŊɩUHwe.�1�S&[�U��I|� CC��Hߡ�����oNz�7��5����S�&�ߙ��Tv���8��qS�q�����7���δ���p��L���C<�X�:� ��1�ˮo3�=��3��>����y�$ڸ��5�l��m����|�e�^�:qI	@W�`m��K�b�~��q��C������ߊ� �^.��;�aai\�T��,��ھ�Fh
:�Z��v#�W}F	�<���F���bw�[7S^�f-CM�0:�ܬ�Q��,c�s37&�g�W�X����.�K��Y�&g�d�zm��\��0A�<D�E�ɏ�"�M� �]�+�v�p|I���EPmD/nX����c���[7����[��l��j0���u�H�>(���]��R׵��˷}L?q&d�K&\q���@�j�Y쎻��E�I�霨.�%r���2��U! �Ӹ��5��Ov- ~��fp,�e�я�|��<��*�_L̕���q)���5+�t�p�8��B|҂>s%ē~��}BEo��g~�Y˫��?!�U���$�MV!�Aޝ6(4'������!�w>�5�)!:�pڝZ�]�Z�+���n[aQ
~#�Ѵڜ�*��܍��X�nj��c�P�)\Q�bT�8�-K��;B�WZ�3ؠo�(_��v��� >�������e�sc�#���i�a��Hc��;�D ��^�5 \��WN%�E)J�0�vg,i�,�����O����,�e�+�Y�!2���н�E�.�X&��AZ�J��i����^%�`q�5����ԮN)5~R�ʷ�{CE�}"+�?@fc�I,,�h����Aa	6�n%�C�j.��L6\����qHМ��9�p���4=f6�,�������c(�U���c^c#�;�2ҡ'�����ϻ�F�G9��قz����M=�J�0
}{-}���ܙ(ҟר|u'���a��uZ�4*���޴�1��xw
��ƐT��4��٫ɮ���砻r��%��G�P�zE>�]OpxVؽ��L���.0jA'����I�����13E��GL�.d<���^I�)��ia�hd���X{K��W��؊�7��F��׻".���Ąi@��.s��9�Eg܁�S�_��3x|��Mz�H��Qv[Qp|����-����}`�@�K�w�X�����~P������ҕ�Q��z�	%���/0S[���_̘�egN��"i�o}e�g����9�W��ӖX��(C�D�@ka��]`�4{�O�����K�Hb++{:��Ӱ#�S$��U\}N/S>���~ԭ��%����ډ�~�>�qf�$Kq��:U0vʴ��ì^�
ﳢ*�3�¬�������L�ŕ�3�P=it�c������ ��/��[�e�O�9E^n,��������b[.Ȇj@��Typ�wU�,�}���Q����
2X#�����90Ⱥٺl�´�T],Վ��(s�/��7�%�AmD�ԉ�pT��<�<ᨻ��K16���}�Ǌ_/0"3�n��[�S��G+
!��rA#�X��I�(���Y�qOD6su�1�0<Ytf��_�PF�;'ٺ�F{LH�
���T�vL!5���[g�o7�	����۫�~������H��@�F8�'8aƄW��ON]�
Z�g��l�����o�'��jP�6��T^k���tr��4\1�Y{D��̜>�5	9���g��ԅ�)R��S\G�[�~��4�,��^y���5Jw��-����p��h���f�r/��k�E��"� cx�4f�c�ulS>����ֶ~��Z�J���w��V��o1�î���~�_:�ʰ_�����H�;�o��?PP�8����V�V���:�φx�n3���R�Ŋ���	�ف.>ӑ� �`���fo����v��m�2�|��3+���D�pfd�Z�yI�xf~��RO�A�ΰ�
���ajC�MǓ�z�hDN�M��ৼ!��0�{Y����Ta��_�=�2$��!����IJ"�>;^kx85�b��Uv��ʓ`F�h�`"���OW��|��g#� %?���_�x8��%9y�����P��2���I�G�R"�tO4���O=d�][nq�ں��P����w��A��j�ϵ<w-q�@�uH�L�>����E��]<�̖U��R@F2?��W���?cS��jI_����X����	K�*ғeU�<IOz��qBK�K�.��v� ��L�[�*"hm@��α�਩r!чw��.[�o^.��.����aH����0�~�W
�?���/m>gv��5��ڿjF�I���"��B^��ƛڎ��$kMq�ճF-�8��3w��s��A���n�n�YK\�l!�����X��>[f��auh:�7 �H�+c����7���{o �mS�R�v�@AB �'��/�A������̦�G5a7���h�V������FPhq��ȋ�}{'�UYZ��^q�k<*߭?Xn,�樖`X��"�5�o`_�0p�o>�����f�u}��Ma5 ��Х����{g���0�r�ȦR�9��3!�Ѵ[��D�Ϭ%z@*��T�O8g'�TX5 ^M 2�y�8���l�!+�gK��V��
-�2w�S�c��U{���K��V��R��~�F6COU:���#BϑB�mE"����)a�X�Y[%��*���Tn���4n���ewd��S��+��I�#V�?gg3�x$?ɿ�y'&,��D��d�g�cz<�J'>U^n?�q8�"���)x+�2��=�UX��6m@���a[�����܅0e+�a�`�}ק�E�%bB�ϥ.D�'S��w$bE�����[b��+\9	���N@�O1�W���z\р@�u�W h4^�B��.J�pR����}I�%E�F�B�o�?����K7>�ld5��psH����� ��.�l�"��n�����b$t�S���3����[V�\���{��������}2��?�,�p��V��i��"|��eD<��e�i�eh�
�Ь�I�w��~t�j�QmR�v"�"��.0#Q/�Hu-�=� +]�tF=�E�e0�M��\��wDn�������T�9	�����ܷT:�4 ݞoٰ�!vW���"����\�!�q��E�7Sb�It�8��a��K�Έ�0̹c��N��>���|k��#˞�cg�}��;��%���俶Wk��.vT�<�g��_�  �Emb�l�S��w)?�{mf�|���x�,���(7�	���?�t��r���*������>���p�.�*�W���i44fS��K4I���Vo#�����������%�si���.�2շ<��ǑfA��If��H�dt�����G���P�fɟT׺z���΋�;�<���?��#�Y�Q�3]����t����f�������4(E�;���]ti�g�綉�#~�B;N�W����iA���Ƴ���F���o�R��ѨH�Bh/�]k.���-Z��|c��{b��뺋���C�pr�Q��<&u�n����v�Q���*�w�!5)O6���;r��ru��3k�x�vՑ������q�� �e��ݓ��,x������B{��%��Li4�\�ݗaH!s�M��W{@��<�1~A���񓞁��c.�e�8M��q�����n'�P"�q��G@��h�H�2ܔHq#�*d��7,�7s�^�S�����������ԓPSϊ^��&��Ȑ��A��ћ�+��2�����������n��X"m��u�2�Պ�^X���kR�����Nܵ�8�H���O�\��C�A@�K�=d���c~HK���9�s��Na���DuJ��6�+��<����.?�"��l�K�d��8�O��d��r
X�v�O�g��[bY�ZK[�4�7��wv��d��jF�xaf����,Q��Q�Y(�#�yB����uK@�VP�a�I_*M,@��|�ـ�p^ᶗfx"�jS3f�0�K�G�I�G}��k�fw��*;� Y����P)��]�>�{:�K� J��P�jQH{"ZmhR �ě�?:�/>0D_�����|�"��4B�!k75�J"�g��6ug�}�������~~д��*t�/6�W [=���rܰ(����]������b��<"�#&���\IQ��>/7
E[�(��w_:5v̗�^����s�a%��I��:$�U�11� T���g�$�*Kj��^��~�r2�"��o�@��C���_�w0q)�� r���T{#@-ma�t��c�H�$Q�Ii�P��	/���|�"�_��;�V	��o�����9R�ȗ%�Mt����C�I&8�Y��T�k�?��I�����BsP���ŒשU�� ��2h`ώ3� ��?`9��%��gY$����P5��3���[�7���wVM��!Yb�t��� ��,��l��R�|/ c� u�X�%.��\�6��2��$�"6a$��� ��y�D��N£��xPJIp�f8���sv��-�;LBcF�`� 
]�'&,�w�菲z~�������A�M�#�x^ç�$-�7������ňԮ@�9|���|�w@݀��u�ޜ�Ӡc�}����ⱀ���f��F �c\�ϣ�{����1�Fi�١I��k��2mk��>E�QVkC���Һ-�ѧD����Ю��İ�{'�P�c�ad(��J�$B��6�3E4LNz��n�k�N��E@K�����&B�+i��5s��/=�"U���W5��<{M��,*��RAs՜ۑ��fn{�^=^;�ur���P�k��f~v��6���=p�_�!$����Ap }�_�.��6�J�_}���fA�\J��c�>oG��
qAr��k��ns�N� �$��Q����1���p� ���pP!������{g(`�B�טjc��JQC}E�tз�[�b�彶ǂ��Mz�M���%�c�H�����\�?��R�-�3���� Hw�{��;��aAG���|"�����LB�-%���P��ӊ�ϯ�� z�h�P)�^��4���7��״�#��Ñ}.��[�T����G��S�J�2����O��2����cVL���	D✓�&����l1 W��Y��T@��￨1�=RЙ*(���BR��j��6�/ D9�p�����v��!<Spu�'���ì�>��h ���'`ٔ�Q<�Y�����2�@�X����ӱ�`���kf"�P��ڭ�#/Q��:���u�7$@��θt���8f-�C�C
��`�mf��)cɣփ�&6���]�(Y��܆R��q�9&U*mU_'Yt+��ͷ:COD"+dE��-��g��%�G��xE*t���}`Sx>W�@��`O�����E�K���u��bc��I�7g/$�|����� ���G��������y'�ry�v�X�=z7�c������aٲ��&e��R�_�Hr�^U�*7�N�,?}�0�V�ö�{-�9_
��@W��>����Ń�@�R�5u7�t����� `�f.���$i�ܬ�t)�A�~V`�r�FE�(;�ճ�E�S�����+-�����AV�F��[�����A��(�z��}L8닀�=�Q�=�߾����X�����^]�h�v���A=}�
7��44��U9X�����7�M *�཯y����K�?Q�H��m�nZ�4�L�I�y-�.�3�`�e�`�'p��Ɉ�P����S�h����*.�6�HU֥+d���W��/�Q�Di�Ϝ�9+�;\�M�f	�Nx��0����xX��~��n�05v��AtLcL��o�2�:�3lZ3Z��9OYUz!r��<�`�:�=�۪D7w��.��g]ԝ`������	Mh�XW]�N�I�x�,�%k'Һy�hn��+Uo�5܅���ՠRi�mN�|��!�\�B#n�9�i��2IBwq�������kS�]䨧��N�g_�",������3��a팠w*ZpPu�ʃʵff5 W7T����`z�"��WѬ/��k*%"{\*<V��˿S�Za+a}'�ͳ;jY�?� Ȅ�/��@!�4����?�Y�s5�j���4�tҌ}��(c�c
N2�X/JQ.ܛ;<	�F�IĎ��`����
�7�|�{�k�J��)F�~ �a.@���:�?�W�P��;󊿙)�C��������n�~�RQ���
��v�p��-m��]v��Gb�vc�`�n�޿���5#'�"���/w��|�_ɚx�t귌�#�k�s:Wj|��A|�Z�fҝ��!�u�V����c��n�\/i�)�cZK ���4�Hqd�e�S�8�?�T��#��/e�\��e��ם����wp��df�T��#��wn�ll��Ro6,�0���V.Mw���4�h$�p'�+�epS�,��co��O�'Y&f0K0���@k��"N�H1��e2�x ��2������
�d���k��_�֍�(�km�+k��h҂Av��E�ps���3.�4|D#_���g}���|�fX�ʳ:��y�J��`�Pj���I"��`���qT��(�+�ɇf�� S��⪯̓҅X���E�y���4L����C�%�z����;��.3y����PH����A���3��MD;ŗ�eY,\EΘH�p�g)Y�Nl�h���b�g���z�h�f#�s����34�f/%3��yCJ���H܎�U�����^��曉��F��˚�d��5)�H[�z�8����D���߷6~24'^-bU��U�7'ۦ9w[��W9W�a5�����|=��g��/O�O��|�Θ��u���۝�����8ܼ�*��{���+��^B؋�j��K�O9�(��.z�]/��!�D�E)��sڮ˲և�X<���G�����hnW��������W�׉�IY�E9�\�n��QR�F��z��~&��Vz��N<T�P43h��$�����1[��7��::�Θc���UDͪ#*F�͜N�A���?���O�ڪ��Qvu[l�2�����\�3��q�RGJ�	f��䰵V���;#�kZb.a�Ч�{���u��0�P���[[�#�����ʘ`+�M�u��5I)����7 ��mö�'vF�=�8���Î��'�����t��+/�yd����ޝvtǭJ)��B�?7� �Ayp��$h��@��H�CG��*C��]տ��շ_t=�m����ֵA������ʟ\��c�
E:�H� ��=�}��}�D�W�~8��<�Vd���-#�Ǩ��"e^��rK�{�Q}^�J<��k�&��c��bld���Ο��c�
��<��ᮣ���V�����z���B����ܚn�zO�8��@xVf�F�����=������`2���/����D �����Q�B��ɲ
��g�L�+b
_ڐ����\�X�V�=ؑYh[�`��B�u8+�Ğ3K�4��N��^Et嘾O!J���T� ���M�-,_��)���c���aM��EvM��e�*M��(���~�|�n��Tt� U+pqe�es'��S��3�������� 9y�"lmh�I�wkf��z������ep1k-r�եS��ֽ��*��X	E�U�K���>��=5��;Js/����?N���/i�·��rcD.��r��ᬹ�J=�k�T��:��2��aEqOWl��W/u��e����K���*��(p|��l���~�h��<0�̌+@.$%���ݖC�U�5�������d��)��r�/�fǭckmNo{۠ˠE=]�>B�C�R_a>�+��u�
�u�����ԧm���P��4�Щu@��,%�iX%	Ζ�H�{�	7K�eD��T�7*�HR��(���跋��o�~9N�b;a�!D*0; H�pݲ��p�IBl��kU�*_�䕚�L-�J�Z?T���{"����턛���\��V*h�l ܱJQd���ͥh�p�օ�ߣި\���ܖek�d�L�w�>cׅO)耧�l}�#a�	�loiվ�:L�Iږ���x�1��h��Ynd�,�]0��<�����4]�4��*�F�u�kgH�r����������R�p������֯L�X{	�ѱ��?��Pg�O��'�,w$<�)3o��v�Y��R0�.s��B~ �o*�UM@g��u׳��Cb[<�T>4 7�����	�ۗ�P�\��k�M7B�fx!0�cb���M�W�����ih��Rg��>[c6��e�h��' @�f�'�<�ʭ&f��*�$�����Y~0@y%SE�G\�*����=cx/�����eT�b5��f�ݗ��f �o:�!	O�s�ˮY'���Jz����xH�O:�'���2��b���Ɛ;�9MB)iP����/Uh)M�p<��� ?�j:�.�[a�y<n
�h|��WUv��{�Gn �\_9�F�zʖ,�7sl"6Y4w�B�Ey��t(��}�"��<ߠ]�ؙ"jiD�8=M��Cۢ�M��s�'{H-׿~�q&��m�L"Q��aҐ�� ������{����̑�*��ME�p���fb��?��8�@*~l�Y��������!���᥅p�}�xx�
>�,�O=�z�B�,;���J#aw� �_ݻ�	�p�� �4�=��MUP�����͜n[_��sX�)����B5���_l�/"��b�S�5��Y�y��w��|:�h������_"�$V?SR��5(G'I�U�c�ʢ�u�t;�bY�jA�����n��`%WJ�L�Pz9�Vf$�i�R3�������<����g��=�: �+�Q�[�C~��u�'���Q�;b���Y��KY��g��|���Ko�9ᶘ�y�*�
+'�V�&���xH��v��0gt���'�K�0J�L�Ǳ�_��s>�C$����y��f�y�* >�S&Np;���8���g��~G�h�>�W�j�'Q�\;!�O�A�^
F��߯�rp:W����@\�?T�`���x!�=Jze�������A�T!Pn;�jͪ�)�HݎG�Z8I���b���s��O�b�=����0��
H���fD�B�7[�Q����I���ز�?��[��i�ԋ���%؋��(�Uh�������M���zH�2�RRu�NӶ���$��e���Kj�ݕ�;w����� ^H�%����/�
xT�Y)Pj�;����B����	x�{<�6����'�DCx/�����Z���#�=�Y(�N�������͕i�(����:��7�O�g��2�.i����f�&��"��t]��]!1��4-QD%(hU�d�(�E�r�Q�	
��#�r�$���}W�Y.b�^S�n�*��B}�k�����4v���Z|r� o����v�V���� �uE��i;cb>�﷡z�H�"�z#b��F�H�v�%|�	�<FD-x��B�J��	z�Y@H�J$�O���G���
P�M^m��&&�W�Rc4����}�>�����mXɹ�����m��!'9�D>}m!�G�̽oK�fZg�CKT���qգw����^	N��yڥ��˓�nⳢ@цꞈ�����ܘ����\ﱦ��~�Y�R7�e�G�@TT&������N����(� ���1]���K�尺�
�w}h5O�壦?rN*�J	�ʤ
�:ӝ<�3�)�����:��
�c ,,���}�s�@�m�#h�^7�2����7!L�߅-A�:�U�Mw,�,��)x���>=pv��l�SyJh&#:x�3�N��@��V|��qY@S�����qA���Ơ�H����M�$`��EJj����:�X�on��$nu�ub~���i�U;���Y�JW���9 o�Wu�-Dk�J�hQ��ᴸ}8byП��%ߔ�Q����m�pl��e14�7�kF������d�k|8���
�M:.:A�9!d��U���{�Z�m�@��l" {[�7Δz?K�{�eA:W�U�����|P6��oq}Q����3��P�B�+�`U���q�����M�W-ZI�޻�4~8����f�tV���;��j��o{�\���O���1�	��o:gΝ��?4�,�o�_�"x�1�(��N�������z���%��l5T�w�� RN�f��%��i�O��EA��;�DJ�c�c�k� �?$��ቼ����7�SƇ�����k�:�.���cD��%��g��P���$��E�Z��V�C��4;���;c�r��Y�=@Ɛ�;��N���	��wYQ����W��Ffsm�a��^�
/�V�mPY�Hb��2"6_��%F�>�0��}�����0�!��A3��4���d�9���O�T%۲]�b��7p6����K&��D�Z�#�$�e���O!���_��XLX�WQ>w�D��cu�����v
�SN�璖)
���!)�cw9��=�#�j��0��u`��Jc�a?*��e�|-�D�jB�:p��$�_�M?vJw��r����E�EL��@��W?�M�;�?O¸�xo�f0�	Q�	���+N��/�X��G&��Ԏ�՝!��6R$y�	mP���ᰂipm��Z:����0i�[�������B�)��~-��ӂܢr�b�)Z����+�?߮3^�g^��)�O0��p��$}�]�㥚�Eݛ�Pb��^s��Y��rzI	�D�퓀���m#F=�4i4�Gp�e��I�@��R�c�D�C����Fխ���#C4�}��>n��(�4h�0��/}�a6�^O�j��Jԭ����ؼ����Tq��ܧ[Ɋ>��GK��q�Nw�_�Dc�������}
Ot�d�C��Y�0�ϻ��`���� �8=sىx�n?m>�k�t	�5Tnؿ_5��+I����Wy�֕C ��6���pp�������c����J��NbVY��BJW���3����/������\4 g���12��\�&�>PW"�#~��E�-aq@�(�4C���:nB�s�)8F%�H[0�Jiv"�.�L�p ����#� ��EuXE�F -a#y=���IE�@�M����c�,����͕Q��C�n��3�U�O"�%+;���`�
������N"�������hm���2����z��<= ��s
�ƥi�w��~�6?���	0�6�4�'��,d���Q}�۾2�hiv�Lsm rH>�oe��Q�k���*����g#��Z���ap(F���}�xff�,���"S��Ҽ�N9->����WK��|���͜3>'R�o�� �<J,���C�H;�)�<d��׿�����P���H�b���gZ߁9�����~���͆�[ ����
 �9>�e�
���*���q斤*&>cȾݷ�~aq^o��F�YD �9�����cs��B�~M @��e�*>ߝ�R �-�'V'G:fɤ�u����0�VA��騉t��wGP7�L�:WU��y,�x!3�D��ۃ��)m�ϳ��i񦧧_�
<�=��A��~Y�.=[�N�A��V��Bp�k�x �r~��De�2�9
���bƽ���L�5À{Ca�|� �g��<6�?bպt�tx�u*X��]<?������+'Xw3����9i7��*m�I��_�qCD��VU|Pn�l�$�0���e=�P�3j��"|y�K֓�v4{t9��'w���/jĘԐ��C�e��f6��K������%<�����|�� �� c�1~Y�K�̴z�YS�9��mW<g���̪�<@�f}a�eJ��ݻIW�z���1����P4�>��5��6&�)j��F.�O����ͻ!4���)�{�K�(g�=�|�-�j�3Y�0Y����G(�ܠy3�KQצ2��� ����O�����oSÂ�����e�0t2����ƙ'��˳Gw+{�"�x�Fd�����n�B3|�ypyMP8B{Րoc훘�L����x���Lq��w4L�*�J�>~��s���e��n�]��+��u7!D�0�E�Q��4"�2������`|�P-���w%�x����	�}�+�&�(�=;c?�
BH�cs&�cH%\{|�&>_?�B�l����7��ǂ�!�6��2���{hM�/� ��BP""�z}��b~�T��X��7t��b2.�s��Z"���bNPʟ�S1��
�{P�;����P�V���}3s1u�d8�c���9��J���y�+�f\w��l��d�	��$��ͧ�d&P��C���M �9u�'3�vb��V��d�V�f(�3e�Fb�ǹa�Od�zC��;��^fI��m@�D
$ &��wj�ʵ-�v�e.��cYC��7U�ds~� �� c������m����+モ�i���Pu]�@�X6�rB7/�d�a*���J��H:��j��ܳ�r��pf��.�fc�S��x��o\ZW[\��\�V������R��C��*<ħ���]�l.Y*=l6��#x��T�7��Etn��C&�4-�F����9�����]i��Bd��Ƌ5	g�]u�[W��G4>�d Q!�Woo�y���).���6�&�����C���A�RX��m1��0H���$^�\9�%���]���h���O�M���|?o>l�09������V��+P�Gb\و͝L�SF��[����^�5��h�9��T�)�}$�J˽`��/�����Rnħ���1m�&������x'�B4�i�*.�X�{��pg�+�������̅]��@��Z�4!���ۣ
0�KS!�Mٳ���!;?y��1/<#�Sgrf���|���8�0ؤ�k�O���ű��AN�Y��@$���0��cbHF���W��W{ץ~�Q$��緒[����9(~�\��5)K�?]�K0w�!��)�,/L HÚ��x�G����8�8�~�b9B�<���ZB�9p۷�y�Ae�8�Lǆl�U"e.Q3Y��X����mi>g��燂?��w>�E��r�:��t�F��Bܿ*�t^F$P�R�9@�� 뾖ί��+�����čJ�,	��=���mu�2�+�~�Ҧ��1"�_��7y��Q���o�b�'�O��x� �\�7 �~o�}O����V�N::���;���X�����&����k3Xl�:�G�D2���8l4����O�:!  ��6�ӵ�%�k6���yY�������vx����x��m��7;xz{(D��e��_-lSD��,��� �'�V��-�fIO�����2��P-nj�p��p�´�M�xkm=X�8*�,a%��EQ>��q_�bB�yQ��uP��S���W ���G�F�����CQk��a�^8jY�1k�A�AQ�P�vs/>���v��7��BG��F#9@���K��H�%��d���~�%�T5���v�o�f�,N�$@hθ`-�M#F��л5#`F%�f;p���in�H�:!�g���)�*�͖[�|��ҋ������U�a!�{.�f�Baj���nG�%��w&M��롤��P|�8�:�"�X�~�J'��WJ��|st{�俦ŘB@5�Ea'*Y����,�e���d^����ӷ�K�D�� y��kJ��Ns��X�֋d��m�J�O�Yl�ۨ��a�{���4��%�A���4�j��/~��ɳ�QV��qX�S-���(���V�z<��r�:�Q%���M�ⵒL�*Q�/��6�
�p<���d
CRx�U���E��߷�o���v�[��H���	dq8o$f3�Ns��?�nh{ L��R|��N�8R�