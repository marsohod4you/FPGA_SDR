��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��։�������7�ь&t����l�e������as��U��p���t��|��=�<�4ХC��-<?_a���}B<�͡��zaRX�oD��I�=�Jz�'���rt
o�G���ֿ}�\���˘�`���P��w ��[*�@�1c��)�,�dP������S���pC�'�y1�n`�Ep�Z��O��M*���lHe���] �fϚIN����~
�&4}����# g,�U��Ȼv�2W|���ƕt7������$ e���j2%����PT�k���uy��~�$��N5��V -�cF�D�
EW<Iy�}	�������l��ݝ+��B��\m�Pn��:�.q�`o2��z�c�C�����Bn�xo� _ �Ǣ�FD^}ZA�S-XP����y�	�Y�R*��Ϗ�� ���R}O:m�� ��9��?1y\�n�͟�k`f檡�A {{�9%���i˰�~Å���ȩ�\�|�S��l�Z& �k�R}��P�ܜ�hX9rV�I��L��������a���-�a���f&=��,�A(��H&(������S�H�J�L%�eM��H�c�9���#	����)�J�z)f�(^�:�ˌ�/�4���}rj��;��\H�E D\A�V[��ص]P%��7��_`]�������E�B7K������0��T�3�/�p��*���ʼ�]�)C�kqs��*����Ö�e�>.I,"bK=Qf�����Ԃ��D��T�gɯ}�ɧ�{c�G[��:�!�
a�L�xA������#��n���ŉ,�v}m�s��#Yc�2�!��ی|��+������ɨӳ�[�E�t�P }�DQi�"�/$�6�,Oυ���t���JR5��sٺ�Ls���2tZ�	셬�u��] �y�H��rYђ2�G9� �p/����;��R�����͔FI�|5����U�ݞ8�a,�xrZ�c�S�2�Փ���i+�$MxN�S�&lfS���wI��e�[�&�����dx~�O���=L;i�����x�f0��IWGL��F�$��2�Q.��ݏ��[&�#��*Ϛ��:��օ��t������E�Omf�� �r�2
�`�aI�ޮz*q�����Ҝ��3�U�H�kGl��YME�T���i�f�4�x��dS�7akB 3�iY{A�h�w��GQ�����X{;��,#�%��"�^X!���~�H�ߌ�˕�>ӯR���v���v��H7b�9ǲ���G4;|���'���*���	K����ɩJy����I���7�Ы��W�M��(	�R&�[^��ka.x�����UR��������\Ab_����i���/)��N�x�{�O�&,�<r����jq��5��a��B���HZx�2�[@��!��n��N>��͏`Ll�@���fWC��ߟ�������o��?"�G�
���o�xJ�f�_O��^������mӘE�~I&"%a�ˍ\'�2�w�*� V��ITXD�=��\���) |sS ?���\��X�}Yp����g�7:th5�q[Ȋ�%ɯH�@藧ѭ%C݉�6C\�k����C�"�GP+��)���/)�'x(J��{�X?TayM���Pi�~�词@p�-�4�5u�G��CY����NvG1��z�(�d?uQ�V��h�.��,X��C3	%�Pܻ�}W���(��ϴd؞sf��+t�������U��(�UA�V�7�C���I��K����hڨ���i����LD�~�S/�x-z���Z)2s�E�=`߸�ׁ�\����y��C`���|}3��W���Z=�[s®I�'�rݷd�$	�?�7KR������e���>�L�Y\���=tkK�q9�2�i��d�#)"4lu��o��ZmC+,p����Sb>�UT|�NpB��AY�Ӝ7N�
�9̀���(ӓW�Fln��'m�ϗu�8a�	֛ t����f�e)(��ox�ލ�"����<�s8`ɐ��"Ԙ��Mqv�+áٖ�Pw-8��(���]ӮR���8Q��-)�vj@P
(�I�ǛgBM���D1=:몢��[4o�ߥcQ�:�ye��E�͒{I�*��!M��EZbj���46V�Pm-X�b�xH��HJ%�)8(1�p9s�zO�O�S#!1h�����r/�$��ɤ ��k���k�hJN�k��r�D��� U�j�1,O�T+Wb���Ϧ�fn������: E|�Tdx��~ͳ6�Nʪ�>#ƒ���)�b�l�ĺ�Wׅ�Ȭް%u�H���F�����Lz�ą���p�����R�x>S�px�������E����9���"l^��b�>��X���#۲�8�:�N�2���E�}N�pk����f�f�`|S���4}����ež�����1��8�*�(���dA⍲�u�F~��٪@��o�%l���Fc����YG>!�iV�|�zv�OIL��&�<lBjF�&���XD�G8*��i��xATq��4�K�V�7/����g��*e>�׍u��"�H?EX~��D���F�	\��7m��.��1���jt-��n�k���:�a��a�U��k�ĈW$a�@�������j�>���:d�"|�YͶ��*^���Sm � L� �򸊥b�����#3?��չ�r�[��\��ʕ��y-뙇��f���[��'ď������`�R��L��U�ݧ��?��O���I�6
�;Ir81gȘ.�-f���x���h�uC1�|�&pd�K.��[%���5��.s������[��,��ď�W��ŴpUN{)Ӫ|�٭	�%�SDn5��\We��`��&�ĕMm��D (2r�Z�g�t��1d�2`�������R9�.Z�����42ٕj��ϥz�Ҟ,�1w�q#��+��^r�H�<z��G]�l&��#���{6kLxB̓�K�'��������:����G�d�٦旾V���ůa�M��j���ȡ~��I�Oi�^��q$�,�R��u��>ċ�O+cW��m��kSם�{�o[Vc����	��������si�*���W~)0����-�}#�#���X��s-�MI	�<�3L��n� ��4�����leho�{U�����#�'D�;�A��D��^�V@ğv��+0��wG�i���:�ϐ��@�9:���i�#�t%���hX:�J���&�D>�|�%�Y',ƛP��+��g�i8�.{���~���dЙB9�d�+�RT���E���W9��_&�
���[EI���'��Tơ]'���Jb��E� �fg�	A��,U��x�ͶU[u"Q�.�������.#C�4w+gi�,�O�S�J��o�Ѓ)z ��7�솳���؀��Z�������$Z���_(}�!����G�u1��N}��t����Y��8���Z�M@̒DP&�VQ�����.����v?�Dr�3¦�u4�H旅�:˅���\�v�l��-q���(*��C+-� ��[}�X!����0{�~��y(?��&K����M^��c���ȵ��b�G�]��(�iq�'�F��x<�@��4U��g���r�u��u��O�����8N5y��XJ<!���h�Sc]6��SC,�C�r��yL�zw��
�c��A����ʺ�R	T�����3^�4��֑[�	����X�aw�ݑF�{FC�E���c�{�º�+N
j��Izj��AS���z�.��.Ԝ����<uƵ���!����K�[#�e{��ȕ)��HŌ���Np��A��T�1�JEH�� �D �T�����P�72�P�%S�b�-�J	sE[��v)�C(����J�k���*;��u� �nf���X_g*��bNW�DpPp�ߩ���(#l��V+���{���AU�Z����>Q�^�
+S�����n�P���^�ch�V�ȯ��'*�w�]�R4-���C]w6H��}m���kz����>�G$m�$�~?ց���Ӱ4�:��D$kbDt��{*k8%���h84�d-��k�>uI'9�\ؖ���
>��R��,]��PW�P�b����à� 3���܏�LT׶όJ0��C�6���d���. S�]18�6���2����N����K��A>�|d�-(5:I��E�8�P�'7��<����='���`�:<��3���w,oR�I�*�x�8Fq���!� ��)H,5u��9s��5�j*��=g�'\�Ѷp��,zNV�)R��M�����}M�����I>4g�&6a�#����9���g����5��$$�F�U�E�]������<����)��g`B4�+U�X ��!;L�j*�p�'��K��`��A����70Ќ%f�]���Z'0��S���w Y��uTϗ��� �ޅh�cS������h]<����h�����	���拖�����@��p��+�np�P�6�������EM/���]�zY�P�	THD��H>򕿚a�=�TG�R�넩���Kw��{���F��4�C�jg)9��g�W�&;���Q�T�nmt�Aw�<��l�K=�Dh������P�Pz'ޗ}���C���"�^��h��=��69�M�U��
H��l���T�R-�*�Jቺz1n*�����ɮ�b���`՝�H��Ր�(��"�Η5'[�k�r;'	��!�O��M�<�����=��i����r�M�_���lC�ؒ��>-W<���r����Ȁ�p��(�FM�R!	д�j���sz�MOJ�����C<坺U0�?;K���&�1�ʩe
o�/ɧ%{�����'0�VV�f���8+�"|B��'��$R�i���/�k��E%'M䶨bV�,�d9]��0��+mg�"}q�/�bx}��G�nkQ4"�4���j������w�1M�r����1六ﺲ�ӸԜZ��g��ȯrrߗ��Ռ*v��Y �'���W(=�QV���Y���/�:��	2q�8�@zFE�$7<q9Y]x	�ʺ����o�s�G�3�i׮�$���w>Rς+̿�v*��)#��N���5ɮ��1��W3��w�=�u���y�EW�@y��� x6��S��`7'�V�/��%�-`w��M�lh��R�j<��K>.�!�{��c��ǭ�hݥv�`ͬ2M/�<ul�8ѯ�gK����>�q(��ݯ[���	L���C3�4�v��O�G[[��C `��qQ��� ��߬��y6�
"�ŜK,ow^o, 4@�t኱=->�#���U/�H4�qy������l������\(Jh�(v1Q�_zՕ���qp$����N{�h@;�[i~e)�x��ݒ�� ��f7��^�����!ͳ<���4D���lam@���^$���^}�Yn���à|�M��M��E�#G>a��-Ag���G���>��Po]{v�z8�Kv�U��D8-xyH@���d^��(e{� � �J�h�y�-#� ��^E3Cn���_¦&����N�K)UJ� *�5tĦ��c-��\'B�H���ɻ$Q�c_��(r���ߐ�9*'.�-W�����N���9F7� JD��>����Պ�3|^�?	}�ܫ=��i���~U��bQN�	��yjX��7ޘ�	K�cd��y@������E�	�Q�.�w�v�U̜�y�G
i~]�
�7"�k昔]�(_�����Cv�V�5t�\\;b�Ӹ5�U<sH��,��Y@|��QDa�!_������#,8x�f>]MM%d���C�R9��&�s|����oYG����g�3�uԝ3@lAh�e���<b�������e����qN��x�I�8W~j��"i��P%�@�h�s�Pr�ЁK��I���3�;��]��E���'�(F4
h�]~�ޭ��%��;<�R�g��"$��:w��0(��wy�(��fa�/K��(�0<��Ɯ���:@�ē����DH��Q�R��6l�|5�B��k7�.�P�� �j�8Xd.5�/l��A�]�E/�y].U�
;Q+���!&��E�}�M����LyZؕB��Fn��AzU����%)�Q ��M?���$	�O((����	��p�PW�P����YK���Q��Tj��PGJ7��"��'zE��jH�sN�
%v���|O��q���~7��*L�v�?$�1�.a����,�#��q��M��~A�y�u������3�P��@h詋v&NW��T�yt��W� ��;�����/��h�w>\5�s�	W��0׋_	ǟ����+����.��V�zޠ���zGR�;(wĦn�=�⍋j�u|�j@>��&d=��L9���u"��u�LA�Ú۵X�9I�� �}�R��y^�_T���Q�/��u!���R��\�q̾�+6KЖ�g7$�ࢼR3����Yo6��6�wۺ���������3��f;��&�M�Λ�dJ�%U��JB������q�/���a�D{H9a!X?��'0p�H�g
�7���1�2��.a4r�$�q�ngZ��Hsʃt��Co�Bqt��d�[vI
ȮW�8��s��O�LY����7Rܼe��HZX?��s�R������G�#��(�F(A�l�d^U�6-8����0�����q��Q�z^�-�h�O%�G�X��������g0IԒ�V9U_�W�����>.��4^��t2q�f��.��
Ϧ�I��q�����i�)�&Q�]�W�?��9 �4����(�
B}W�Ft��mq������Eu*T`w��$��|5J� 1�h��L1/-C�Qݱ�!'���oo����&|�%,{��1_�dzC[�m3�"O�v�z}g���O��E�T�χbT�[�j��J��O��f���O���l�O��SlӞ� %�jG��p��׏�1@����F�\~��a�f��ּj���U�0ܒP1�y^��cK6����>456��z&�g-d�y� XT�ka$�;��P24��\6��G��҂�ۣ����.�Wk���9s�[(���j�30��#)��^�NX��a?�p7��@���	��[$��tV��j�E��O9;/�Χ�R�u�w�ָ֕�{V��U���ʂ�Ez�P�{%�);�Bz��&��]i]˕9$��!�MX��������F�wyl�.Aֳ*��6�L��ڏ��3t�%�k+�->�z]�)��*`/��uK�>gg�v$�N