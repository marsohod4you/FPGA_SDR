��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+ھ`��+�$�v���NF��a�ᎻE��u{~Y�B|&��ky�t� 3'{\�L�*t ��ˇm�[@�(6�����?U8p��n�6�
�0��2��v5��	x8�\�^K'.gFh6ʟ{���2�<�#�u��3�U,fI���Qх����
% �B,a�(>����������k`�N���S�ec��T�z1��ܣ�?⬃X��H�*�п�}��t��1��o|Vr�NF���S�֪!�=��Eb#�O-~A�x��p��B�_ߗ��7*8c�<1v����&�'+�n辰��g;&T1�c�K��9�1\�s����iH��YΜ�����y,S ���0�a7i��j���
�QQg.ܘe{
#0pb<c��!q�#/����<�����!|�O����Ѫ.t�U����4�_hc�ų�]����A�73��̏�����P��d�K>�c���S8�/����E���x�`j3�P`�%֞9q��UX��:����������//�J��[ML7iu�f����X"��S�#�su���n��	Q�jZ"�##��
+Q�m�L��KZkt�D�CR������Ъe�_��M�����`��YK:��)*�D\�z�̖րC�E}>�3��}�h�~͊�L��*�g˞�s��a��ʺ ��ɂa=�m�-�@��a�r��b)�T�q�w��p*rB]�� v�Y�t�yך�u�V���O�X)��?��1�C�K!�'�2X�p�(��ȳ�5�f��8�����:ZR��5Uѭm��;����>1�C,�k[��Է�'�����l>��<�������>q������~��C͍��K8��!�Z��.)b����Z ���� ��@�v"|M�%A�Uh�BeDƎ�&��R�J7X�F'�a�XFqo�n�w��s���845��'k���f�3��V��|2-γ�ܩ!"�X���ݞck���p�f�B���Uڟ��[� S;�:�2#�E��xW�o�����=���Ώ�:���A�������!R�� �@N
�	�#W@���T�)����	N��X�X�B�����
3:`�q@k{'�
�����*�[N���AZB�@4<}L�B(�cݯ�n�+��m���+dA�e7�C'�(�����`�lК��:Ά�t�f��Fو�[�����1z俬��S�R@�d�������B��>��Rڧ4^��Xu�#}���B]���ƿ�zh�zap���Y�譙k�"�<�ߊtE?;��������:R�eK�*�%����oX�B�_���`��ř2a1�����J"
b����
�͘�Ʒ�(�M���s��A��%���"�p����Ϛ̤�3�-�"�x���Q�ln� �a�1bC50aƽ�D�u��,�,Ȍ��L.����D�R�B�3x��B~<{��L0Be�f!��_���&w��n�Rʩ�/�:�&,C5������p����,��*蕭"�w-r��$���pl��fe �!�W�R��N"�.e>(�I���*
����HR���J�*?L߼�|b��e�C#����m�@�f�Vk8�c�P��CaW�/�͇�d�\�5Rt��>���:�t�%S�u�(�'7����د �Z1�S��yC��	�;ru�PIt ��G
�Ȇ�#H|�l�՗�z�`������׏�K�~Zݨ�2"�A-i�};���W
TD:����jek)�c�q�E�k��?���"��w����^������#�Qf�I������ �H`�ҳ��V�N�O��ڔl�����n6��e�0����)�G��p6.<U��Bׅ�96�1�m9��}�C�pQ�D��[]�.򄫏���~�o�c��c?�w_����HRB����F�!�b�,T�8E��뭒ӛ���H�K�����!��?�OwP�i��f�Ǝ�>��S�G1�me�oS��W���V	����֢=�9��A��_�����hy���߬��r�~&���p6�+��tU���;},�kyiv��`5ĭZ�H���qK��^	ݚ�.��AW�x5�/R;[7�?9�f�[ۈ�����Ǔ�����Ԑ�{�S���HwQ:�x֕Ԓ��,���f,uz7h
�A��~����ej���X��s/������G �j0)=f|x� �C�H�q��x6�?���[A�-�FNW)�U�E��3���Z����;A�[���j�mm�\�w�Tg�'�7v$��dڔ2�֯:��R���\G�Q�߅����K7��K�q9���l��#�\H�1�[�nhe�}��/J}N��3�c��*��~��\�0��u��o�,}!>���@g?k7]qQe�x�2.m]��}�3��#��L�]���^��ލ�p�N��N�C�@�T��Rgb}�]l�t+�ez�X�:�a�X�aGD!E2�j��x?>�<�7,3�]��s��5 �$t!׮⃃v��R��A%�?�G�����U�+Z�l� ����@o�w'^	�c��U��H�YA���#ҁ�-�2P�u�NmV=oɯ1�/S�C�~��$���ʤp��w��n����}�>U� �vHrC#�i�.�z�Q�-e�ot�q���BgCH�e�z�:��
l����;�]}�H_m�t�-U9`$ 8_)���ਓ�ֿe�gTv��2�4 e.o�S�����
{����cG!��o����'��~)_w�3Y��K%m�0ϥ�x:0jy|﫷;��}:EP�6���gV��\�
_�rK+$�62��T}/�	)���b��������S:'����4��1p���^�-�:%I�?���>�7�g
G4�,Bm�����<׃8�m�q����`��6z��g�Q���-<F��*���0��h(W�ϓ��@�"�^�l��ډ�H��CBq<�����D��'%�W�P9����V�˶�)8�����n����4b.���X5���~'���0�EՂ�'��)gҨy	�:J�WQ�N��D`�J��y/'�q��2��(rQ&6��f��7��@��,��9d�s�R�H`��5�3�7�l}�a��Q0��ۓ�>�({@X�s'�v�(�����@�L8�i�L��V����-��Y��`�rr�4d��Q��xC�.$����J�Ԇ�{��;Ov��WWg�4�>�k�1�8��0�9Pt%�/\p�6F��'��
�W�΃�д��ˋϬ<ƭD��!��c��Z�
�'>%�F�\��ʶCp���tj���v��
��j���&�C��������)J�)ʐ�mK��i�B/������o`�^ �Mc��K�2u����ڞ0d�{�����z�\i�Y��r�KU�
��k�i��n%(Id-�<�����g2�.i�|Jw�,?<�H��$���Ŏ���u�L��A�t0�A��VQ��I.�aP�b�d�mEl����B��4�5.����	Vx�6�j|	�YJG�= ?h��B�`#x n(��V�;#]o����	'��Ux��<�E��O�D��ӅL�:2y}o�g�w+�8>��C��Q�v���6���=� >wT�1����í6ڔ�|$#8�j�R�觀Rӝ,2ajp�)uy\L3�c�X�-fޓ��:��˾L�)�7	��!g���1�s���#Oڐ��\���HU�/�O/�.�����p�(|�6��G��Jd?F��nTx��g��#B��&�p;�0��= �ja���^��d���\c۫��FM�>��Yb�XNo�f��F7��wN�2yf��l�(�n����'%��{���7�?z4���`��49�$�ƅ�m>-�_��i(T�=WL2Ϗ���y8�8�U�u�@�A�i��i�<ٲ�*� ��m�j:r�D-��&�^�S*Y�@�-S��*V?��5����sH�ij���iZ���kZ}P�\"[i�*G@�f�pU���"�m�=��`W�.�$Cu�d�PY���W��Ɲ������������LF�LG)�ք<��U������rôx����W*ѻ�jQ�^"��6�;����r
��Fm��� ����UiIX�b+j�;]VAm��@���R��$@����U��9�����^�"�(�����o�s��/�)o1���l�~�v"c��ϝ�����z��?I��o�Z]�ơ��I�E88�)���wA-�R�t����	�<u��Q��P�St�n�?�`��n��o��W���j:~0�����:}`���(r��k%#���"Qbc�c  �+����\w�Z�!`���4G�$)��h@��@�~S_�̫�\��%�V���_���!�X�s?T^Py[����=�(��i��
ܠ��\��9���������: d5����H
��Mđ�u��[S;g�EK�f�p�04�烞q�"h�����wz��Yl�x9�ʈ�h�'�:�Rr��T����?ޕغ���?��o����V�haĜ��HR�650y�2	�����C��\r��Y��� $�۵��*�#���fgh"�n兼7�#Y�a�Z2u�!C�F~�'�T:Zz�nm.��[e��4'7I���z� �6�*�(��б�-˕K��B�=�^��<.�����Z+V�b������Y�s�b�e�����w���]�5+��y���q�A�,Em>5O/��@�ah��Jr+����0��dʷ��`���m�`[Ry� Xؒ%"����o����k�N*h�L*w�D.
��SN%�}��$M^���:����?^&��v�h}t���ʹ׻F8y�gC�)��n���S��9e�����"M�T<�0Q���_0�ϧzxw���]}Ϥ��[F�j��#��	�"E^j ��]�{�b�ܜU]xI���� �H��k���ՌzK#F�ѪD~d�wG��$]���0e�{DF�~�0����+1�1d���{��8��(JpQ����n���<,���4�v�#8�D�������7�&ka�@3�׀�I����x�(GXXʮ`�+�7ȟOL��+G�!&
���U��P��t���l1}�mK�?#'|]��_�"��C#^�l�Q���%g��y��'�����3�K�)��s� �%�fa�� ���a��\i��{�*�+��{�e*k�\\{�Cq���fN�����ɵ��oi��K������B��8wO�㞅z��{���9:J��~X�B��<z�<O�qU���"�O��'���Z`���J2�
/9-zPy�]s�gk�U�1S��ͨ"�!�T:s[���=0���u���i�>%�k:��j��h��'�a�Q�?��H��]x�o\����:�G:�{#͵E�f14�ޟX,r��M"�l�Uk��]<�`B�"���?=�(�����1Lk-(K7;��7�h����&.�H�(�ค��bIh��s!�'��{���.J�{�׋�e�o:�Ӗwһ+Q�fL��5��1S�oam8�y'p�j��Ѽ��f�v�i)�����wI*'i���?������{������)4����o�Ad}�c(N�ڧ��!��#T���'Z���c
�v��&���b�Q��vR�[�Y��/A��B�H�[P��r��X�����ڷ��'�t�ΣSmHY^S|��l�b�
揶��PƤ2� q@+e��W��A�22�'�����X3�#xڥQ#c�\������"���$m�;�r}���	F�>�>;
#a,��r�+�i��ZR/ņ
p-0�F���;\��-G�2���̅� �6���6������o0���ͿB�(d��Y��L&����|�i���//?�I��J>���S��A8��2 ��@� ��ڸ7�����]�e7;�F$3ؙ7��7HTwFIA��4(� ��š�82��Vm����no��dՑ
�2&_��T<�5�E�#��mH�D��A��Ԟ	���UI*�<C_�i4��V�S�).h=n�W�Xx��s�ifS������ �L�����~?�f�Bu�������舐�B�Hf��u�^rf�L`�U[�␕��=��	�=�Y�q	����~(}J��/lʫ!�vֲ���������d����*&KS����� �!˛���}B�6t�8�N��	�10��Ob2�U�U�7בN�Q
��l��>���l޷hF�Z��F�U������[��$�sE?�c Ň$'5h�:��E��j���5+(H�h�ds�3��^��^��O��~.W���f��IG��p���+����4˯1�}2(�^]�f�^(�p1� �鵍��/��e>���E-�'�.G��