��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K���e���c5�B�s3!S��s\:=][�*��7���ƃ!K�Q���ݠ��۲}ͩ�<�>��>+�J��ph�m@ҧC���9*/�5���2]R��L3�(��}����0�$��O�-���"8E��>�<�.:+�6�X�u����p��MdJ�/��։z�Ցł�U�`�4{t���� 퀾���B����6=f�1�l��xSa��S�[�x����,i����;)_d(�l`x�p��\J	#�}�T�M��H4>�7��؁|��r��/5楆 ��衡P��YS�7A֢}�n��#�B9� W3#'~�3;�M�cs^��9��5�����2�u��2�{K�V�W�iuR��`8��r�ٽPE-r��8�10�N��[��?��V�Z5U��j�gЏ�/��r�v�������DԆ!�xJ~�yƑ
=�dޔ��Y���rS���1�[@X5�A9Lr	)l�g����>��c�X ��	C���=���	OYv'CA�.�ۇ���-�d�]I��Pj��qk�	N[<>�]����;��,��]��J��JrT�}1pOC��w M�9��M��P���E��jk���ɍʿ�;��w-4ze�͍;8�K> �hM��&�����p�	�1$�H/��$4m^ѕ-�/���7{n�U#�#�t���x��m5b�1Ef_��a������k<w�m��.p^ݙ���q?���4�LS��?�̫C]���Q�B8ޔ[�pXa�}��w/v�� �x��[��ؼ�L�P�?5��Y�2��ɩ�1�2im�_3��·� ����Z�����y�`o�Vڭ�wf���-���p��6<��Ңl�Y��U0�e�r֊*aƜQ�w"D�B�<����K�4�}?>C�gw��)��ǯ.��*4KҍUA����#Ցb})s?;��'��Si����`�=�кH�ki�!hk�X��^y��j���}��t4X0�P�X<�~6�������(B��LQƢ��o"�_�,�4m�wu�����Lj�J��꩹::�F> ��2$�����z���u�r��\4�^�
�Ro����qT9o��<^����A��c�ea����~�I�@>p���Z��贲��R�n�Q��pY�	m��ҕ�5
~r���J34T֒��h������*T���GЎ�
}a�_����������~��\Y���e-'j}���`��J����f��܅�kld
~)��C����g�P�B��s��g"У�e�9֌H���<K@�!\Jy��ͱ�YS\�����4#����Hm�9��g)�?M��'�)��e�
��"n��W*Q��tT��r'���ƞ&����vώS��&%�,��5P�sS�G�M k`�����b���#��2!�j�㼶;սN\vRrܼk1[�G��L�ҫ��i��yQR����v�Kz�A��}�Lh2�z:��[�p�.i!bX�����B��ơ����=\A��8����)1(�b����1�^g�йz;v$�^��w�D ��~�@.+)�Q���X0�:�>#{�Ε,�`񌥅���ţ�>V!*h� �jq��3�F/{�#3����CԬ�<Cx\�
���_�	�Fy�x���FK�� *T�����R򹡨��N
�^��g,E
a�[{���+�	(1p�1*
D��/y��"iĥ����7���m�ʷ�_�R,Ӂ�f0��W��j\��N��C���
�/q�h�p����ui�M��fR�{)T),��| ����U�5O;���fp}�=���f�T:%,�bS��)!�I'q��V�q�S�Y%d^�&�{����*s�A�IDK��-_Ӽ�6XX"��_9יs��-�a���b���*z�IM�P���/ꟑ���K
��b�lEf�Mq��j}�dp�ɑ�=���f�vt���Y�) ��56Z����do.�뿬BFH3�4�Q+�5���R�[le㐌��땨�xB��� ��~Q�?T��oO1�V@0����R*� �ʶ�o������ٝllx�E)�ڱ\��dшϨ��8$~�mf�x�r|�����i,l��"��b;���r�M�'E�z�T"� ����JR�*�幙�i���B�����<	��@,V��.�l�g;ZM	�;��w)'����"�Z�Ci|oɋ�v��[O�;���K��jJu����`X<��{�U���@��#?:�R�n�������칮сĝ�p]2����]̼��I�%�ou�~�,����� ��!�"�����z���_�-
)fw�[�����3gI�� m
�#��x�N�z�<�a?lz�"����-׈�_�pF�b+���a�`"{�M�
7�>в��=���yL	�E7���i5#��Nm��؎{��"y�ʗ��ZM�9أ��/4z�K7�ax`��3���ރx�;[��!���\c�ɟg}��T���"��Tb�FP�*u�� �ھɧ��n��7�W�
���eD��g@HC�L�E��K�՚<\�#��W�Q����/9h�:(L	�9�M�ֻ���Q+�,�����u>m�:g>�(>��Wу�����漯ib�ʱ�s�O������f�tT|a�f\� Z[���Wi���rY��&��q�c�}��|K�xk��w�����MBs� t��������5�^�[��[;r��L��LU<�������񑺋:�z��hm�]6I	�G=݀��u1"]V�~䚩ȧ�@�.��z����p��wBE0"3���rG��(q�27T$��
��0r�o�=�dv�mu����J���E��~S��Nh5��R�rۀx\�!�+B�3U�tF|���[�'h5w���d)���BI�:A�>P�~��v�<,>OH@�c���*��B���}?���Z(�rs�ۼ��J�a_ͦp�`��I>$~���j��q���3��tpˊq[Tq��;
]�|r��h�b%S�v,�olx��Q�O��Bv��w1黁h+�4�^%�g�����ntd�0d�;��L���7������*
�?��˅xp�����&/��@!��1$Q��a�a�U��yۼ�D�⊲�x6:�T�K��yW�{s�Xi��T��j��k8�W'�g�N*Q�b!Ծ���s�n	�7p�������m`��3��V	��D�(k¿����M�VF��)���:{;�}�G�3u�/+eU�K�,�4����8�Gd{7�eTJD�����-g=t"�޲�o6��,�9�9(�E/�f_��Sw�o�ֻUA�^e��Sp6��4��W�+'����G�w{s�RTdb<��^�wJ0:ъ����x�!�v�'�jD���><����'X�m��V:/5ޗ�q�՟0FD-��F�Ҏ��-��Nю����
pm#�E�ѿC6��@���
�VO&@��N����t.��R �1�a ^�����:cKz��U�AC��^�N�p?�4�.Pb�ł�v��Ee7ވ���%45�l�,����ӃO���/.���0��CG���r@��M�����a��qL��Ρ�e[�P��j�{ci�g�|��i� �+�1P䵃���LF�|z�#dC�e��	�>fP��FT&�6�up��v�7��m���ە�I	� �#�-�����6�*=L$�����;h�
�!�������0��٭g/�~k�QV̀�l�#�A�`p c�B�+m����c�u?]�L�I7�dm�ʛ�
�x�؟{�Ǒ��=T�X��i��M�Z��.��̯�3���L��KY�A Oq��E�U�д��t�?�?z�TFs�en*K��U��0�����)�4r��B��/�O�^��N����uT���6���,���|�Q7�����#5#�?;�(��r�W�F��X���^��ja�V�Y^��bE�`+D&�_�`	�֪��-���A��c�����r�)��J���+�y7;��Wlϰ=��%����$�J��,<�#{p
=q��i|s�͵X~��Au�Y�x�;��g�����+=+�,(��:�ᩀ*o@u	e�ӊ �h�O�é7�mr�?pֿ6��Q�J/�UV<�	j�2M2�sr�7!�����?�mT&��s��}W�7����n�QR|{�Ti�mP�w3�5[��E��K�1���Ra>�,�����2w���;/܃������L�+(TY;�T�xF��~���YQ�Հ���lT[ �Y==�daQ���p��G���j1�T:�A��
�yr�^�꨽Ғ��C<��/�]���Z�G��/N�s�|�'?���+�LU�a(���;��������.`�dc���+[5����5��$���H��j�����7�!�ԘU 2��Ѫgl�7�J�S�ԋj	Ă��_\$vE�h�^��F�� z��K���.2zw GP3wp�&�7�=$h�-����]CJ��>j���D}5�e��ϞgJr.r���1�8_΁�9���&�^kDb�ˉ�"��"��+�c��'�/-����Oj�V-ö���ֻ�!&���e^�����d<���+i�8 �Aҵ���dV]}ϕ�k��������+J��s�}�c�����]8`�����@�R/=�yg\����Ȧ�R|���Q�����1�^}�t	Gܷ0��HG���x�a�$5�
6�4O�Z�,k���J|���� ���&�����ڇhW`�����?U15�?�O�-B�0a]�4��8�0��VӗZ�Z��\���vuxo�NB5S8���Y�a���a*ᘋ��	��K;�^��  4������g��BlȮv|�m�`�N�V-@��fm���q�"� M\�J�������.F���Cm^AV���;����Q�O�C2�y��VYCz�2_9A&tzci?=X�d�d���?Wƴ�ꋿz뾞�F�|k�{o7���܏,�[���mk����ۀ�A�Ƣt�	����V�|�<��K�h{3�^�k3KD>�(:$6�u*��������(����v%w
\&LQ��b%�s�J\�Y�
&pW��}�����K��?��ž������x�����I=��8�O*��� 3=n<�>�,&�y��<-2�_��g�;���x`k��mQ��%9%'"�
�
HL.*/���d��\)f�T�	����w ��4�(J��ޖ'9��U}J�e�h������E����]:#�:_�甠�i�3�;��>��]᠕�NIO
�/�z���M��0�
��	�>/<~Ju�%ۀ�q���A?��:}[���b�#w��������������9��a
ַhE�P�U�_��Ld�Fr�4F?
���$:Fo8A�g3ġ-6k�����KBPހT�u)n�x�lF���d��g���I���<��J0�OΠ8WUF~�Y����!���iP�>��5�9�9���l�����9��q+eW�y`�[�aA�]
���m��k5&����K����/�=ے3:�EC@��k������*�!�_Z��"��	i&���#��4|E��[�ڨlӤ$yt��ט�Vϝ�"��To��;��%~���]��9��|9Vn������u�Z�E�c�2�]2i�#��h��a�U�CĜ4��VY�k��J�n]��|�sH���K�s����x��%K�+Z@h.�ڽ�yc��О�[��/]L}M������'�=eվ��y]�z	��t�z�nb�7#EO��:��g:,���\�β��;���0u�%�t���I�w���e��ۘ9l�ۘb�0�v1l	er,!�-��2��u��b�w�3�Z`I�85!b����D���v��?�a�m#R�&�ks���>�{���{:Yu��e9����-�W�,p��ަYS��O���rp�Aw����+�A����0���w��Â�s�5*԰}�`~�C����j�eC�.��Q�j��L��$
�#K ��O�^LNk�X�1�:�s�T�N�|�����a�ؤ����vu��֎�b�1V����wD�J���"�ʡ�w~l_�[|��H��"���d�m1��[��>�JE�őZ�{X�/���J��:�F_��U9�-�(м�<T����r�9�<�2�$yڹ1.����BP���]�h�J�j��Fg ���"|�� ���U��0�4h���I�����YR҂ͯ��^�k�EB���s���46�l��Vb�Ș`/\��9=Ϙ=B>�͏1ŜF���P�o<7.�0���2V_�/k�	ڛ�j�_��mU����"�o~��9���� �,	�09���.��!YJ:� �CB�(M��n�,Y�1�*���G�'V��"��^~����\c}^��1�U��[������b�/Pi�v�g��$~�ʢ:7�Jn"Υ6���3/K�����h�-K�W)���3Σ�'��/�&��3��[��㱍.ud[O��~(���^��.&��T��k56�s;O]2W��@<�����/���pX�Ki����^�1*;� �"m��i�`���b�2��'�3[�O��&��V���G%�Lg���S*����B��x4u�#N��VP%.�"<��+�n�X㾷v�K���-���p��ۦ����̑��O��2:�v�0��0J&�T?����5g��GJ�ī\�����[)E�^sr���+��D���kp
�0�#VR�`�.<���>4} �7��m�t:�X̒�=c��F7ߗ�$�o��[�J���{�����E4N!#ɹ�f7m!��y�S6�P��*Gኝ׿{Q*k�இ��`Z�yf>����sK�u"w#U�HD_r��Fl���� [���=V���8� #aR�����!I��lJ���K���t�����醥C%ov(#�*�PqT��|/i��/� ʴ]��j��H�̣�]�U�|*������<��X.�c��K�j�B�F�1Rl=v�L���������T\'|��q�����b���ן�6A�,a����?$Љ��@��3`a��WIy���iH�_�Z� E��^O0����S���N� ��X�:��2	��k���"��2-A�Yk���LW�pi{�w�$�~�R;��jQ�P��b�W�v�ї��PUFy���z_"m�Ѣ$�E���8.��Si�JBU�P�K�7$�]����Z07��[��C~��ꉏ=kۖ��vE�e�iw��{�K䓟��,Mj������7��J����t�l�J��4_)�*�� c�/��fN���~�&�<#�1��� �g5�,uj簴�g�_����Lt�҄!�?C�͔��f
��e㽘�W���`��۵Qp�k2�Q=�X&U�C�oz�� Q�M�X�qU�����F;o�I,&-uq�j��e^��� ��Psk'��d0�+h��Sr	8
*6�- �ӅT�7�C� Ynr��N�*��J��'F��X�`ge�ash��,�YT�J:�#1���ai�|^U��9�h2e)!���e���D0N!s�:��Q+�E��F�$̐�z���9��!�����ų%��>�/Ɍ�_��d����aoe��妒+�I�"˲0P�1�9����q�c� b\W#��N�qI����J��� �}�i:I/䀙1��#����q�2���x�E�?��v;sXnj��{���Ru��tH%������0'�3#�3�>��t��`l�):
�p��FO���]Eg���-�!�����6`��@T[uB�v�^*^�TYq�H?#̪r�\�5���Ȧ;��������G8�$���]t��]�y]y�R�REX���?ߜ(TD*`���!|�����<R�T�t����2�O��RA}�ʚǶ'LR���N�����_�o$b�_D�xz�/ y�a�ӳ�.�пFcZ�8�>�� �L]4Q��G�E����@�@[�l����]�ꑰ�5f3⨚��N��ڗEKFO�-\HIO��J���~�"�Gi�=��'A��u;Ąw�`(���k��~�Ԉ�qX����oh���k�<�qA�����^u�H��9��,/=���S�-�L�L��U�8�?4lK�O�i�.j��+�0��W?kV�5�c���,��X�H���3��@j<N눔�Esk��ҳ�i\R�H�덆]e��8�l�7�v�Vz�:�<��������j���4��3lţ�$�4�ޘ�7hA_��N0e`�,.9�(Mw�I��9�Lf(��a�p��*�-I7��ޓ,�� �D({D�E��a6�j���
R���P��l�`����boqu�i��-�!��e�E�Rf��x*�Xf�P�B`��%�X��6��\^�]� �/qx�r�Q8d��Cː��x��|��#�N������G-SL(x�]E�� o|���2X�6�c5�,�e�	���?%O�;��]��[��N�Kq�I����3�9�ĸ��﷙�����1p�$�B�u�l�c;��8g�f�9�E.۰ne�_����>�����#��&��Y &-�$��n��,)����0�fñO��#�Wk/J���D���|��w��<�L����'YQ/d�����G��]�_z;E���g�J�oRr^V=�q���hf���Y9�#��q������Z�F���8�����T�k�a3j�~󰎗�f"3�j�˯{�D����
��|u�ǄJ�th�aO声�J�c5yD���X��+]�K�ء��>ţη�=g�U��7Y{I��
]):�btH��V�y�: b�[4U�+J��6JjU���i���4�n@�xnt�&���pd+�!�\�~��y(�{��x�f��>}�RlF�ŖY��g���,�Ϋ��E��י�X(�)�A���D)W�,>�%�>a��� E�R���o�6X.��3k�HrAџ�>���n�NJ?�&��S*#wr�	��Q����5�q�Zr�n���pB���:���)}4���H�I�:�Z���>Kѧ���z$�C���h�ʥk��Y<��r�gc7z�%:��|!�^c?���1N!!�K��5g���O}W�I\QC�|?u���1e�6Ԛ@��|�)�A��y�d��Z�	��w�[:�BD��~Ca����~��NL�QN��Yin
�w^i�SS=]����{���r���ڮ\�<�*�������]ɿ#K�l���)�J��Z�=�dy����i���i��V�u��7zU5��5{�2Ea]^3�P�P���J��&'�«���=������Y#b�B�Hr�9�(^IS��[)s�f�,,���yK,�a�� �>+̝K&>��;�h�֘��	c�N����w��58�=>�����Q�~�N��&���_[y,�u)G��J�|or�׼x��S9_��(�_�a�3�-���,�K'���v��v��e�U�������\�j iOo��f6:#���F�
�ݕL*�5"���@ĕj$i"�Y��]��m�^Icկ)#6%_6"���ݎZ���*̉Yh/�i�'κ���<	j�Qbf��]w�C�cf�Ig�n��⦟x��4�-�xo�s	'��J��ש%��0մ2:��Z���i��j$Ƚ��Xˡ�	8՘��DFò+�U�I�ܶB�F��h�
˫3�5��R+	P!bQaȉ~�+D<���l>d�� ہ�;9��aH��S{XUDnI&��#Bt����3�Z���th{oci��?f@Rn��c^�N8U�K/�;��
���us���+�G��J�#�D~�-ޟ(��8a��5���7���j]>'�X�*��ύ�;Muk;�ϻ�Q�h3��4�h*�Q�<wGC�0b�[C�Z���u�Z�W����)NS_�ٲ�z� (ή�%�@ҋ�;��6_�6��^�g�L{��^���Ѯ��`�}��hك�yaU��Kᏽ�8�	�s����8��Z�6*k}QK�.�h�ᾷ��2��w:!h/�F"�,z����0���e�0��T�q�ʻ�ה�v=���v�F��>�	���B���0�Q����U9SB���	NTB���?T���fQ�ϔ4z�'�=e����;MjE�	�����ξ�._Y�`��G�tv�[`;1}����N4{��v��\���PEi�]P'S���cmd���%4�/!�y���#�������v�<C�Qh#@6�g�_�ݖG����Ƥ%��a��ED�Q�3ھWU~�ZL�X|E�f
�Q���4^�]+����^c	��D3�7 �Gѧ[�	��E⹒�j|[��VG�{A?w����]`��%t:wR����c���"C��^#ާ����	eaXi"�J�/Ϟ��x��i����h���Vɉ��)���7�w.^OS<���~�#]�����Ɉ����?�)�XJ�/��hd�;��4�ػ�	D����ju�o�ʱ���{��z�X�Y�źv~9���Jc� K�Ҽ��?��{Pb �UM�8F%UY:9�m���w����^�Y�L7�αWk��3�x^H���'� �(��f�x�;|Wt�g��
�R�4n�y�����;�8D�j�_(2�2�FM�Sm���9�#�#�T���5x�X�9��|���O[�f4�Ś7TPD_?�T>*z ��v��c؊�� �%l��>܄:Z{�j�kl;W"*�*��1���/+鼯���A8-�兠1Cډ��WG���l��dZ�|u�O��R��|lb�1V�����%��$+!���~*�U�G�@]?]�6f�|.��:��Ey..�?\X+��p��J���S����q�2ț�tD��[c�J*���)�މ�?D�d�h�OY�4i��|��Y��TӺoj��c"���_v������cz�xg�.�ɒ'~7���5c�&V�[S�|�Ll���%Zy�&�w�oՃ�1����ԕ��z�H��$V�ej�������\����_*��e͕�yDi���T`���9Z���@�\Z�!6���u�py=�܊�`$��nC��eѿ	�tKGUc���x}
V��^u_�=��3n�P�K�(�`����t*�7q�����x������s�]�f���a6��"ε0�F/+��gV�
m�4{�./Ņ�jپ7js�f��vm�ӳ��m¢�?y���S�64�9߱�T݋��0�ym��M"F,Eߠ F>	$?��f��TV��F�ӌ-9����Y�C�T�k�S����'���A�\��&X�-?�V����JBLK�d�//P��ǿ�J��LeFW�W�gW�d�b]}ߠÛi��&3���[�AT�����*�8����>s��B�r�t/�6O��e�쪋"�)�i