��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ���7�dA=��p�Ȥw썀S����?8g�*��'G�>�����=�1>�b�1z�v�'y��)��{�2.��R_��]JLJ�D/|왒^�V�u�B�Qp9[^6}�	��7����M������g�]��/3ٌ�K���к���f�GM��׎^<�8d:��k�����Ef���q���1Z;r�Z�%/8��H������ՎA��j'�Y����떴a^��	.o�ޡ�b�>Ƽ<o�W����U��=��i�%��K�\r� �|!օ�Nj���#�Vaiޑ.�"����,�=& ����|-�;�\|O��w�&j����1oP�6@����}TE_㏆�f4�캮�M�p������J��6��;�kT�2a�_�_��N%���'��A���NNaT���,#���+?��'��p�b�Yl싂
���S[�!��e���:f̓�7��;��9�%���6Æ�=�asv�،�X��p�e<��+L�[�q���]͠��Qlߌ����o,*\���7��X���Y�K$�����+>����ę�*��O���T�w�����uٲ����'z2�����E&��^�Wa6p?)O=��o����N츆;�
B~,�\�/\<n�c������Q���so״&�'��`�OXa'"��3&�&4B�b�;ZQ�� �Ē�0�.a~ה��ͳʩ�b�V��z�C'M	b��W;uէ#PH�,��ɏ���Ǧ�v����>�4FD���i���i*��h:��6|��n_-�eJ���G��I��W���pc1A]�����N4�:�����u���ļ��EgF[�6{�EĮ��;����$�!q����_N_�,_r�� �>�f�tesZyY�j�^���>���ku`���zs��P�{ʝB)ѕx�hm��nJk�P�p���}#!-���u���Ǽ��҉��x����]hF�		 �M,��g`���!���*����=7������ �qHO��X�>w�$8O�qU����8��Gns.�;�_���9�T�����z?k~E��כ�&���M�dlUV��Ǥi�s����Q@#�<iF��!m�%Ig�~�X��5�{�������C���kA�7|"�X�(�Zc�x��Q����J�߾���ß��[�0�ׁ�M
���;5黩�{�.�$������0�8��fGAX�\k]<:i�_�l��޽��z�|��.����&��@O�HK�s�g�C��t��N��{K�uxr������s���P-��j;ў��� ���T[l�*�SlC������c䊎�J}v+*PՕ�M�Iԓ��|����<��̩AJ��
|��u�R�d���h-8xz����:���� ��Msԏ��J�Ͻ�C����U<�<"�:M|4\�uyȷt�7"xN�L�	Гj;�fA�������3X*��4���h���"�q��D���^�^P��&\M��dv0�t�r�wB�f�_i�\�i�����y��ӕ��6k?&u��o"O�1���=��1n�����O����BI��\Z��pXMqy+;Y�q{��M�����f���4Q!��8⬥bS�UP���q�,�e Y�C�����cs"��<s-(�����$~Ql�~�L�����U~��3����\�}���Y�94
oW�b$f��IH �d��)�K1�k� �z�묅�c�.i�l�,a��l��ژ'�u�|q����dF�zKJ������@b�C�����Rd�0#a]���jc��������k��t,��j�3�١�NsUi�y�"/�|�S3"Zp(�Z�������I2cڝ]:��G�U��k�P��Lm��SYl.��:�;��M���2��޸,�i�W�����lv�1��>'�T%r��T��.$�S���T%XQM�_PD�q��Q�c�� `$�Hz�����bgb�t�$�'�[n�X���j��1Ҕ��T���1`
mjHr|Py@��;��W���8;	��� �ؾT�e��`���UpG��M��#��Ao�����̠�*�׃�*�;�2ؔ�|�������j�
�	��������P��ŜxPnW� m/K�9���?�k�n�FM쏓zVt=�E��d���V���{�PЗ+�
>2��>�G����8 ����h��tt�kЂ�����.9���S��2	>+�`T�yq���6�cR���/LאRt	0�[k��/��"W�]�ZŚ�,�u*�k~�XF��C
H�Y{���1_�c��t6n�:�Ư���݁���}P�:���瀊T!�N��
�7!��-P^�=F�{I25w8��i�|����NKg�!8yw�\e0��j��4v9<$zli���g��9�x"���a���~��V��.��W�I�F�f�qxiA���RW�3%_#���D^�3�!�����a���r+#�Ϲcm`B�����$�f���
��4OV�Ζg�Ǝ�z�G,�V$8����)`�\I��X�V���`�\Tʻ�9��߇/6b3e�[4I4t�TJDz-��ہ�̀�=I��Dh�QA�.C�y쪐����I��(?���>tm>��;��_��#p�0C�^�+}<��CBAC�W"�K���|c� ��,���M�)�X�1�p+*��Vs���H����g��er��hG�;D٪������m{�{}t��!�h��~�'��~��]׆�jiU�rB�#D�� 쵽9��X$����
?�ߑO��`u�wu��*���/N�.���>*GwY���iJL��Ξ	�����JQJ�)uPf���d2��^�r��]��'�m)8PW�~Zמ�h����Mv������!^�e�}D�`��ΰ��8>W�j�6E��QT�MB���B�-�
���<��������{��&�v��i�B��M���5�Q��*���}�G�ʫY���$U�����gZ;hN���j�غ�!	dy+>B���J��&ܿb]5�����4�= �>�q�n۵�x�ڐ�3�[���~G��57P���Z��X��O0��e�F�����[?�SM��PS�����F��P��0�zk7ŝ��j!��泾N�J�+Sw�F������3�݉����x���,c�}��ɑ�&���Hu�	�F�INuN!��v�=���⑂���CS�]#���Kr�L�~�� �h����uE/�!�P�-7���<����D�+L���2�ཏQvuK��kt!���a��]�d�G��L��6���t,�q5"B�skꔙ��ٍ�m1�V픗p���{C���N�����	G�#.+L#(X{����gP��u�(R��F]eBm��z".�+*s�*�r�J_�R�~s9���u��b��"4�Es�ñ]�-]�ǚ^��U	3��V<R�'"�q�7+���Jy�)���Wz?�kC".���Sy�п����:��ć!p�":5���8,� �Q"���;�Y��c�s��4,Fq�
��#��7�Glw����� {���S�3�4`�R������n�d�ꨉ.�5�a9`0�h�{��B��f�B�� I��U���t��P��^e��WD��#^N�C����~r�-���!���,.J`Â������شn��b����`&x����Ә�\<�h��-(�1I<\�P;�"�.�4�93���Κ�-m,?�Rҽ�!9��$���w�.�f�^1&�!´�S!h9�%0�	m����}�qsg@��#I({��;i�I�kh�����Ks���i����צ��St?���.SV!eN� �㒕�}Ze�ȸ�N�>�C�z9(�Q�����mMl.hֱ84 :�����떧��Ҏ�·u*��z"x����֖���S����#S�:8��Z�)�|b�Nl���}�f�NՔB�Fhdm� ���L��CZ�.�翗Qu5%�t*�`�.�Y��{��ːERq,1"���H5���(�䓅���d�X�p6��t�z�Ʃ:0�F�O<}������s1sX��Z�;ģ�t�yؑ�o-�~{�d�����߇�;���=��H��i�Xo+�r�V*ִ�)�B��l�Y���y�" P\����P(u��hk�BQ�$���	/+OvI�N��g
�j)"�V��UB�����¸��oe@	���L�:�M��H�f���i030/�Q�ʸ�����X�f��1Ԏ�kԦ�1��,� ��lM@��|�����^��ˈw�$-}қzGDC���K锍IX�I�Ʊ��1�	pZ�)�%�#-a�	�0���Ay,>Α��!��?�@�<נ��%��O���F�*UQ�����s����yE�^��6{��D �N��]��,�w�UN���6ZH\{Q����E.��S��$K�۴Ȟ�LA5����wW߲�e�՛"-�x �b:W;�0�T��d���O��j�{t�KUF�q_Q˦�"�5K؎���jm���uX�I�E͵����ו��aV�ړ�/AN�X#��B=(�DX�~�4���iR�T����C�`��HP�Q|^�GN~��@�	��0Uu���Dl��IKy%w*�Y^:8�p�����i����Ϋ�Ͽ�I�@��/�T[%����B����vʶ�񃠟L��L]+ڬ�	�v`k^�؄_.���a��Gl��?����$ȡ��DGoݖ)��o� Zk(��q�t��cY^�$Ppr%k=����,�j�n�B|�Р~��*KP�!�>{/�@��t�s���U=4X�WO�O�'���m׳o�y�EqE,�iz�+�[v=�� �1v
;��B�����y!4�+�;���@��Sl��? \��@��	��d*H2:�"	�(��/�'�S�*r�n�K�hg�/��fwG?��*<���0��J/u<Q,����A���8�42�;���O�g�"��N��E%Q�gg`�Fʉ��n��b��
|( �4�ý3���ޮ&�'�ƨ���i���8���&ڦ/��_��v#^��#ȃf��k*\Ĥ��7�]�+d-hl��둛k��:���e��O��|[�%�_K2c�I�y=z�t�c1�*�-�/����6�,�!�
[��*AI��C�ܿx�d�c��דF�u<mI����Ҝ܎�
�6�k�j��R��U ]�6#Ҿ'�������h!j�O�LRʷ9�p������a��v�p�/:���d�a�q&��=j�>�ЋX/χgy�OG%jɦ���|�DI�J���6PfC.�����j���%Qx���<� F��%eo�K����0߁LH:�HCm4M;n���=�|-����7c����Uz��2x\��]ւ��O�s7��y,��i�����?=5{�����P)�}�#������u� 6g��v0A��z����n�9�v�v���/ϩ!�J��8.`�^<��mL�,�š��91��\�����j���λFliܩܙ�	�#4����`��X���{�gO�RW%m���7�w9�Z�Q�_����-�������ǝ�S����ާ n��i�M|c��2GgU��s:��\�ކ�K�K����Ng��8!;�1�:Uu(!S)�aA�;���s�z]Ӭ���Ju)/��YMoc�c�J��t��I ��5���W�	��#��b*,�¨�3G�(97��F������������y�r��y��~���kD���0���F�>��ع �t
�r�P�l'?V���`��};=�J���!�7�ϟ0l���F'�$q$�+@L��ql�#��ZהԪ����l��(F2��C�j1g��f���ٜӐ%#s��*m(aB	g��Q��]l9\�ti�����
��g����R#���&���(�R`�_�AU��~y��jBHz���눇��-��@�P�r�(:���������)%��W��s-�=>`�R���H���K�KE��4VeB��X�j��7�N^�����pLX��Y��� ����Q��	Q��Z4W�����L"9ѐd���-��ا�?b�X&�6�����V��_��ړe�l�۹����M�g�ˢ�t��2i�Z�cG��,��M(,]���.G-x�0хe
PCR�%j�����gi*&�t���r|�a]��j@�3=����Y�Sa����+�$���U�-'����ޔ�G�\k��E+���2�
�a+��ϳ⑀g���xߛK�y~lV74�%MO+(]�q(�0!��~4��\�~��!u\e�p�E o������_�0n]^w8��Xf�s���9�h��W�.H`�G�\�!��v�[r��ptu�� 9_�j�c�jo�Yͪb!#R;��n�a�)�ǨM�y�)�v�4¶yڠ=7���Bŧ�	�\��K a˷+ ���	��*�� ;|F}�j��/��ޔ��R
wMu�� �(Z{�$-׃O)����깐�.^c&�y?�����h�A� ��$3Ԩ^�b��^���]�`Lu�<��	m�wx��G\8�bRnk�USy��
n�c�K믠3��$��(&i�Ϸ2�]�:�����E�'��gց*R=�R�Mq}u�i���+�8J3���i'��r�U��&�<��UƙB+��`��𭾆����k�����Έ@�f��N��x�7�8ڒ�*l`�� ��8Í�Rٰ�_���L�Dy*Ie=#W�EI ?~eȡ��V��"��i zj1k��K:�/�@�b��m�DẢ^+�j�� ��Em^��f
�3kW3�4����¨��q9֣4��o�1�o�:���j���?�a��`�͟ *�^�x �&
B�WP/C
{t�Ȣ� r��%gK���ỗ�N�)�K ��4�`~��uy*]�3�ӫ@0�� �ߐ��ʚ�py�����Z�N�?���>�Q�CwR;��3��}�~*�W�oyk`�L�cϲ!�Xm�_�E�%��o WS��M{�XM��(�1ę��[�T�l��rv�8M� �0�j��}?
"�M�~p�u�r�,�=�Y�8��_%m\�QQ��>T^D��?��^ �Y��N���k��H�"����Bs��j���:�	{�2d�7%������~��/� ���lB*|����A�,R;��/�&����Λ�}2�a\ ��ig�M��1���� b�W;D��i�ou�%B��>Ѹ~ u��z�{����5�Ɓ��R�E�o]�8�廇|�X�f�3�Q���o5�� �U��=y"�1����!�����ô�ys�U�{��r鳎z]���}�V��cuD3gП~M�4����F�eEt�a����\i2���ZT�`aͽ�vFvr��K$#�Q�k6ײhl���ٜ稭���ب2���ʻ�f;��*$��T�y���@Ry���h0A�F+����=��A0�R�Y툽MF4:�m`5|͎6��Gb�3p���߀�q��<!��X��*�����4S��Xn/�%��@J�������eT�D�����k�g%۞9����0IX�����MO��$��x_��f�\V�ܻle�an�b!_��0���ٵ<��)5T�Mt:�s�PWq��Bɚ�ɳ�;��ߋ�KP��������w�����B� 2�!��Ӏ�O���W�O��';$�ۯ�.�i%�lφ���Y�4����]�f�R�8�jR�H4�ם�X���8T�M�ŝb�:
V�.Ub�Z�c)Cf�r��+k��nJ�?�i�B5���������@�UV�Qg�b��$�* MM����p.!���wX<Aa�&DǭDa�z���EQ>ȃB���~8�j�·���1$���9��A`�M*L&��eOSx����=���<{��,imF}aL���tyh_0.AcU�N8`0��G?�O�8�����&�H�e�QL����޵:]�bȱq����#�J�q��6�Գ�{��A��i�^K ������[�S��zӇ��u�=�;�͊��^4O= �?�8��$�ѷ�?���]��3}�+'ߜ�=�|MoH��s-:#7}�de�LDM��e�[h�G�-抏��췶�C����)
{�Ȥ�O�|QE�!��c��w�뉑��{��;x*��^��ORv%c�3�e!��+�tVh!�� D���s���n�U�+	��8q���?[ʞfb]�^�c|@M"FpQ;�g�3.֗����s�W)0:�n@��r�c�ݾ��8M�yܱ�U>� R�n���'s�"�PӶ|6Ç�Q�Sѡ"T��M�������㌲5�'A�uR�z^�@������a�������>���C�մ�$�����@A�9S8�e�,��j�ݖ�GN���e	nb�Y��u�8=M�[6�_HbS'8 аp��_-Hw�D��08�š*���-[a��O�[]E�A&/#ݱ�x&����P���<����|��Qqѣ8n ě}�X�z�ν8S|�tqڟ\ٵx�U��M{*�,�EuG�CȽ�k���n��:���k�o�\r	F_xP���MC̝´�:H�<|H�mc����� gx<�M^�����j�Eu%��x�� �9�$.�̣�P�/ Vm�B���W4&�����{���XW�vl�R���ωWYz����s���t�L ��qɆ�:���rH��@;U6h�Sj)%��X�����=�73���e?ZJ9t����R3|�d���"�S�������\@Qp�C��G�7�����*�i��ldȕ��[���2��L.�=q�v�͂y�s��?j�R3�u4��:�2�<���b�K��*"�v�����k�2����&V{ܯ��$)������<O��@)��62���R��"sXhx����WAdB)̙���m,�D>�B��� ƀ�6B���mh�dE]T��0��"�8$[�r��޳�\<��|����"D�Oz��z��A���-�UA��(��|?�6AQ(��;��;U����T^��`dRf�+�G��Jbc��S)�C�3ס��ډ,�&��
=@�R,|�l��ϓ����֣B��gD�DLR�љ��@hl���a�
r�N�';��j>I��ث��T�"2�r?�C�������te����<{�Se,.�m���S(M�TF��K( ��*��i�1/_��~+��$Ĝ��h�uۢ����+��r�,I@
�p��{h9�.��\X̳��[J�'�&{���	c+2"-�t���4Xa�(b�Lk��iZ�0jp�
?��F�<�A��ZS�z�L9*��鬍�Au1H��c̯��-cL��b���7�S`W,����ֱ9?lѓf���	��2�+���i���s�!�LՁ`��CȰ�fD��k��F��E]Շu-�Z��)�a��� h^DM�Y2\m2����f��J	Q�>A��({be���v�#��5���F]�yu��9*+6�}��=�8̥=G����6I���uK��(�6�/e��վ��pv�/D�`M�Ƕܭ`c�aU1Q
���@~lӀ
�@�bPK��ǝ:����V3���ǝ��`�	xcçڦN�����N2��w4��0�T"I�떁�g0���냞� 	� 9�f!�6nwn��d]&�]�򍫴F�v�� �if�s�AT+�@~]� ��5�F�����g�f�7(:B��F�߽�𒽇��B5)�ؑ��i!�4�J����ޟY�?v�@f"����r;��,-ldY���aB��2&�j���[�PD-Ryj
)|jg�0�dG콕��?�6�+�5^�%�\�`��?.���?Hu��gGh]FHAIa
҉�]?�׍V_֤�(>M�`�~�t�e�GfT�G��X�*d6#H��	��+��i�ԓl�PmǷ<��b��ɕ$k�{�XEu_�B����Tm��4��Fڦz��:F'���m�}�	'�xKb!�9{�1/�3^iHь�����a���nt��;��z̖�$�w��?�B�?�闽i�z��-5�Ɏ�S�0<74��L�ꂦ��ue&�.�h4Ti>��P�d�Bu�u����,��i�"PRg�2CR�e�V��T֫�\^��_}ZT�7�X4�����.Xۻ�y�(,#k�x��5]-�)�#1_&�B�ｉb��Z=t�_���W~����3>�S���J	#��m���w�γ	?�Z)�y�#ylF���dӁR�cq�&ݫ}��@)��~�(�?��pA�R�Lpx�R�}�8ˠ�S&�|ی�ΎQ�zޣ����
���{[�y=Ed�_�бz�g�����U>E�r� )$T�P�����Kہ��#=� ^��8^V. f��|';��y�#�<k��Q�3m�)� F�;D�
�Gf��ڷl �8t�D�X%�����aO'ō������씇
�����͈����&����m��ݡ������T?�Nvs�L���Aoh��7'5��:��W�V�3��H,��9-m��͗lؠ��|�����(�5H�<�����s�AyՂÙ��"�h��؟��쫅 ��^�5���r��p>��-�>�i؋�X��+�=��6ѿ�t~�+|@��C�b����[�y�s��=�Vq���p����Eг����ØP���G����{Dg��8�V�Ȫ9�(,�dl��_�7єr���3��!�v'1��i|��O8<�i:�jj>� �ɩ�P4f����k�)M�䡵䊾spҢ�ߍ���4ڲ�؉�&�q��������a����+��4���\�;�<"���<S��g�xV��uVd��vk���X��7�0�w^��}m�m�nq�!y��}
OF�d���d����t\��F*i|�tJZ�b=F��Ӈ�v����~K���\�R��ͯ7�gX�[��E}��I���]��#lr���N
q�!a��G��Uq�~��+��Pj�9KWq\�:D���l�����i�3�a0ݭ�m<X�2�7��zްE���_�JK��N4��f�ei�����_�Z�#�F�G�����v�P%�=���R�;^����0�R��<�Tg#�DK�