��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>� 0�ʪ�E|�$�c���~��K����`-*�Z"�3�ג4�J|^��k��R�b5�huͮ�*r�q���U$��X����WB�+�	@��%�M+��54����j�V���u����a5m"��G���Ac�B��.��Ȍ�z���yAu�Ф�nzPO=M8���@5"y���GP�,�f���91�iH�9�xsh��>g�+��K!q/E���UåcUO�>���&��������k����"s��;0������u�g�8��
4g]C���5�Ãj}�*�>]�
��濅K8�*��n��#|.�p�{�Pw�rYx?�"#�P�Y��r����������S���ɵ�_h��AR1͚3�ɂ�5v��87��ty�U��G|�MQl��/OV8�=Ѿ�_�7h���-���x��BQ�\��H��vܯ3�+��?j1�[��Ô �"af5���Ņ���F����52ƔЄ����\k��BD��:=���t��g䕍��	�N|ȜK���^�%2QP@�(� � A/��}��F�:�Q���<iU�3�`@�"���I��P�D		�n����c0�5F@/wd&(��Cz�����
u�6UIV5��������b�nUkyu)�x6� ���A��?8�}_��Q�+&�y�J-1_�ռ[%UB3���4Q��|`ƈ����(� �#&���SlYز�}�' 7�+iH��\�]��d-��'�{��2���L��@(�u��U�����N��dK�G��i;$/$�@;o��	���e�"b���<p�tz"��M��,�%��[XJ1�D����9㊘f�e��ZLP�U6������䝖�د������:�R�֐!��zL�S�Cӟl+����0��)���!˙Š:`�GV�1��3%*��w�ԦwX�4p�n�>J8a��P��ʒ#Y���]���{���g���y�LV��p���fҿ=�M��l�ty^�F��*�����w2�4�cQ`5^�l];��L����0��}�x'�'�55_)���j'�'�q�p��𤾵����y�3[��Ҡ�����f��6�Tv�O�q�(����4	,e��E�(y/���Ơy���5f��U��HȠ�V}�f��L�GK>�!)�2n� �,��zǻ\Y��gUb�O'����Sdq�� �7���o�F*D7�����P���F��[%�V����2xfa	~_-��#n]xb^(` ��_wȅ牬�e%jh�4�@��6"��-ɺ��]yےE?Y�����p@],ڴ���}��/����\�F��u��U�5 �M��ư%N)�ঢ়�++~�� ��X��ۉj�<�ߙQ�a��vTBh��uG���?<h��n,3E��rRU!��e)�v�P��@��@6�^.7v4��&�y�!��N�M�f@�:�&�y���R/������Xҳm�����.��tjC�P�Om�(���l/��1<m?iO����U�~��Gjܦ� �{aOci.^G��!PY��
�oQ�_��!���z����S���8������ <��%-e��f/sse�,��"�)}�["�A��t���J�����pCqsj�ڲ�����nj�<%{� ���;��	<��3F&f:⏾%��q8e�SeA�S#�jD4/����\�=^'�=3Jh��\w�"p܉�X���?%�]���,We]V��E��w�~�r����{���3�o�B=�f�������z���!K
`�'L�B�&"���������������ZS���# p�"�8�V��g,�B���R̺��q�Ǐ��t� r���ݛ�7��@}����v���9�� �A�s�d^k1��j>B�t�.ӵ@9�ƌ�1R�2P��U�;��n��=��m�'0h�j��ܴ�+����Q]+6	[��%잢J�D��Y�n�B��g��q�Yٴ��3�xPDʬ���&F���7.�@��F�sęF�^�~+<ZM��J`��9V�) z��:Gy �-MdB%ݯ��U?�u%^�����G��5�賸��g���
{ ��^s��b�8��$��
��=���Nb#������d6�2���D�Ή�a����o"F
��!�*�r ���=�s!������ՋbސnGZ�����Q~t��Y���]Ƿ���%��
��k 7~����[��&Җ���l��p+������7�i�v�b�e)�wG��x�!r�aPc�`��n4��Y�F�'�u����	-o����`�G��)��vJ)�\AE_��(`�g�����Qh���vV�qmXm~ed�蒳���,%��B�$4�&��QX�}�,%I�(s�;�j���E5_0���Vz��,��U���b\d.vm������Q��V���95�L�'�u��R�YCƯ�E�}�L�U8�+��A^#����͠fh&��~5睗X~����h��Q�t�;H�G�����D)��ya�ˍ)�>Ȍf�D3Іd%ں)JS��;�X���`ޱjQϏ�����57��kt
94nM�B�Rv���v�v?���O���Sg�d�X�.tt���Y��yo\�^�wP�6迉�s��qM�8t\�����(�Ɠ��iΩ��+>o_���]R��ʑc;��K�]s@��m>�1��k���@�����Z��k���tj�TG����w	�%�)�N�%�fnǍOqX��{��A��gv�~Ob�)�W@��b.Moj�ad�'��K0��n蘃��/�go�����(#��d���P��+!��Fk	���y��?`����|,�X���Cc��XV��-�n'�����}�tX+�ĸ��D���̚�4�{��Xa��r�ٶ 6w�
˲]�5T���2*R���7�� cwQ`�q�S�xV ���n��Sa@��y.����%�������:H�eb�H�y�2U�6G��/���oj�պ9Ch�u��n1���|�Qox��=xpO�&���������#Hq�Y7���"I�������
�2S}Z�m�/h˺rs�Q������@A���
7�o�vp�2����[�E���@1

�'y��M�Z���R���$
c� �L{���h�9���Yx�cI?&?��:pĮ�6j�~�#9]�QD9��Ί)�A�[ٶEd{�J�*��ʗ�<�8�Qjwb��&����x9
`g���c��˅_��O\8<Y��&���E�S0��;�M�`[����D����hH��v£()U��,C�ԣ��P�r��ڍ��m�I�-ms��w�C�*S���*F���o�(ش�ݵ �V��YIQ.��]�N];�Ԟ(1