��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���{F߶��&��ހ�.U�>{}��}v�S'����ʢpn1aQ�R��4&Pt3��O�	��i.#id�&�1����Z�����)D4J�=T���#�ZwYa,qy�����u�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0�&@�����h�9�-[�xa�A���D�t"s�
�fh1 �0B�mFL�S~���)������a��UX\�q
�h�Z@��9�]��X�-�W"���T�3<�w9m��n�25
;T�4|A�ip�4�ge��Q^p�iU������T�k�	$ٓH���!��Y]�"Y��Mkt��c��Ch�&�, ��Tɢ%6�(���Ipi�C�ɀ9�Kn$@t�=�Sr�zMcy���td��d��T���b$p@�Ds�����j&�p���%c��>I)�����X$!9�xܮ��+_���a�ڷ�X?@]N��� E��^R�M��RG;��T��I+��Ɂ���Yq��:�]����zVխ/�ޟ&¾�^��)}d`��nw����z�4�x%�LӉ�$�{2[{w��L}�&O<m��'J��Jq ؑ�U���_����句ѓ���g>Bu~�8�;Ne�$Q��pތ=m�l�š$���������O7?v�SrBQ�;�m,�.�����H�(��Ƿ*�m��%M*���S�	WU�|=qt���G��Cg2��E4�Q����#m���K�@ �\�Y,�v�P��(ɺ{Od,���R�UˊHد� #����I6Q-϶1�j�Z���*����*����]1n5�l�YT���wR��f"�d"�Ɖ��9o�b6W���A��)�����ܼ�뇭�}l+��TO��Qn��f'���U�їj�_P���=��vg��a\C��y��^k}pE�(�:{��醄boW��>'~�x�f1�4�y���'M��X/ee�Ο3�`u+�C�7	m~pPi��lu������PjVx
w�<)t;�'/-�=�s�S|Y�u�	|�ͻ���;�*&Y�3]>���� ��?y�@T��A'
)"�<�Z��Q�s�2��a$y�R�jH|�~�*���Mn��$�U�W�<��ۇi`oH[5ɸ���S[���I�ac��n��E��c?��#�����%�L�G!+m&$��������t���{����m�>|.�f�8ّ�S�6ز.�P,�qd��T5�U��m&kB��;�/�q����C��K�,�5��P����?eoۓ�?�� ��Vv�z�'!eφ_UW��+��(K�%s{f�X��q�s��8)��(��cE����a6]c�Zvi��$!J�� Z��T�ҷl�`�����'�������"yHZ,޴�6��'dɷ85;_���[�w�__ߦ�
-mY*w.��]aX8Xx�P���ogv�t��^,p��d_`�}�s�e^�M9�B͏���[԰kZ�T���u���C<�f��Y��=G]-�drԏjC��W��&���.qu��g	���&G@�:���4�;o/SܙT�'=�y�qئ��#]_�
��|ؠ��A��)�z�h��Ө=��`\'|F~6J%4΋8 .����:J盯�mh�@�U��V-x̹�������p.[;�m�1(��i�j��G��+��9������&?j�����z��*c7�r��a�ǈ����!��5���k��^x��a�8h��t �\�޹���1l	H��9��Z� mE��W�� �I�6�{��c�1Z	�����Ө{�3�wҮXqL�Z]N�ğ_E�x�jļ���a�r�uC��cp��R� �-GvV�r���4C��u�\0��j�n�pMZ�r�9i0Se�����W懸/� �y0q�����dp��4J`���cP�ໃ�F+M:$z��1�=�u���|�U�Eރ��*�¢@�]�	)r&͛C�V�k�q�. ,�׫��T1cYx�f��`��C1~`��?#?9a��9c`��}�J�K��T���i��G��!��ϼq��!г�n����(Gx>���Ѳe]L�]� Y�`� �z�T�FUX���좈|��T⯓��g�����*��<횜/0�fl�/@B��ђ��m�B����-��pqv�#<|�hS�k_J�<f{u��R�^ß���y��8 '���\{X����1�p��������w�?���_�c���o�8ޠ�7_I����3�̖j���C��<�̮q��nQ�'�M���a����L�p5;��Q�����K��
|n�Ų�������_�p����*ҷsӅ��B-���Nn�F`N+oE�]�}��h���3��f�ij5����Cʕ
���T��Iie(�4Q�Ŷ_�����k����[
�zIl_�����&�zW�^���R��	�\���<���(���}6;L��┮w�:,��P��l�SMx��5�טx���Ŏ[Rvb���<�3��&��CY�`��:�� MH�O������8��R8y!�(4pg�O�4�i,eU��ٰF{�����Va�/�ͤ!Ř��M�rP$VX���OB-d�Z�`"��~-�A��{�Kҷ�"x�#��k�w�;j!�À��Ӧ��&2Gc�j�}'u�!!��ttKY2o��L�	������|_�&D�uS�uIՕ����� �55�`�
}������db�w$���a��+buq�u`��z(��X�P�:DZ�MZV%Q��^9J#oܮw ����5`�n��6yU¼]\�ե)�@��:c�0���qR/�#.������>ZlS3�e��2����[!ޅ�1���q���ɻ�
̴�O�O�8���YC��j���I'2|91�_���i���;�gv���{�֩��R��e�����!J��8+5\�e�[j_�0�[7�r,� ����� �C�`8�,�e系����\�y����5���z�v�Z`X�A��Ŏ��oCu9gu+��v�<�5��i��@�-)a	xAr*��(*9q`ƹc�Y��ʹ����I�r�3�F2���w��F�� *���U��o­{v�`ۤ��G8�e�`K�E	�� ���g3��tl�5Y��c!�X��>G�_�Y[��>gq���l�Y��P��jcq�F��bn��=���\8}K�ܲp��Q�wu�|H(g�;�b��h>m�Q����c��ᐰ%�T�G}���g�l2s���9���$O�~)���	}F�r����M/������6�m�ju���u��:mnBRe�ՑW�n�{Q����֯ĬI��:���t5ʳ�e���~�CՌ��`�Y3"�p"�͵Gܶp�,�:fU�ژ>�|�đDfa�%z�L0�Y�caĒ�F��i�=Z��S_ԈN��)c�g��(���\Qm]�#(�?�ڨi`ϕ�j>N��˼��AF���|�P��a}����$��g��*�%�!������Y�	U:��U]�،�n�l���?ab?���M���N�?����G��p�;{{y����V�V"r�C������%ɔ�G�xb���[Z���LNV�5��w
��K�fD�$3ȅj��.^Ω� r�y�6 �VηO?G!E��a�@'���t�.�{��'b5zL��=� ݽ�9�;�
���U�7�lG ��,h��[�<��!��C�r�ҩ��h4H_���7Gc�Z:ژ��Ս+���m��`�L&�ҟ^Q�K� ��(k&S��adT],��ּ\�e��9{|�Y��i����1��(l.~Di?L|#���� 0�M]5N������c��
C"��o���t^<'�㎟�c�g��-�׳x�C5��$�6���ã~I�x�x�n #�tf��d�J�����g��l��~�smV��Pl�pC�ˑ/p�8���Û%2�(6K[��M�^�����\�zyz CS�A�hF*���GY7�d"W�����Rp�:�����',M�j��%Wm܆��X��0Z�&��PLz3��qr)ۊj4����b�T%%=���Ȍ��s�=c����2�AT	�Y%����^�b'i}�b ��4�;7�G�Y�5��hI�=1��<��H1��X�ʞy��e��n��cճ�%���+���e����M�����(�=����ɖ:�1w�j?��~1/#��0���8���c���0�Vɰ~Ȯ~B
�%`=�n�Wi[�u�n5P� =$�D�Y�88&��+�0M�6L�[E�5�sfS���a�L(����sOq����͈�a%��p���M�0�AK�s�[�D���/� ���%�*QƼT*�0V��۫&���[[}��D���3Hg�=X�ڢy8��Gm�����+r*�C�(�RrE�LE�Z ���kyT��;�U Q���Ќ�e�<�E��XH�yF�b6N��&k�m�z*��`��1mt�1i�+���h��=%Yg%[�<�@�T@
��d��˗B�]Ů�[v���<RX������qa�M�J*����9J�_�<�u��1$����#?5m��K��r��qik�$��Cg/�Ϋ[~���aᦥ�]2=���D�y�6����1��6����aY���5��(���04��|=�}��y���qO���6���?a�:��}�}��/(%����MKn� R�h��~���>�2$1�{�Ć!���N�����HFbAYB� x<wY i@�.�7GY5��:�9��pt-�,���>Ɣ��j�ö���~Lv���vt�ZzJ7 Ȯ�y�;�R0g}s]UqLב�j N�� ��b���;/�8t���Z����@!���*3�Q���֮vtA�a�p	��U��6���O�c4d8sl��}X?"���\q>�~��OS�G>Z�z�&>}�F�NH�j�|�l"
��%%��@�p�����OIfS�%����ΐ���)�|��,Yco��מY�= �h��b���c�[)��h������GET���΋�Ic�Zj���"�`Y����UG��v+�}A�^���R��`��S2�h3��"�}xF2�_���He.�h�6��S,����^X�4HfW��ګE���Yf���_�Jٗ�KQ�F7��=WUK�Sfj��$���ki/.��[2WP����}�Y���M�G��פ9k��U3�$-��=nj���u����s�i��������d�M���7٥�b���ī,�`���5�fDXN���?6�׀�ړJS<ތS��y�aj�$df����N���	��1�6>��@p��琨1ֲ<Łc�m�%,�����~�l�za���~3_�A�^j{���+����V����F�tN��)�I+��p56m)�ճd�j@o�
�qm1���ڎ�i'����p`e��l���`X���_�?����A�t���L� �1�@���v:��h���g���v"�>F$�h��)� �2J:	�Pnv�J�j��
��o���U �ڌ��=d]�MU���l�ܸ��t��eҘٌ�q�ĿD�F����n���e���'�9x}�EWWkK��>���~�&�[c�(�@�E�tk]��dj��F	AONY��1T��S���iU�q��O@�:�f��� �/*8Ux`N���E�e�y,�@ ����
6@�M�o�uR������=Ӛ�}
�:d�Y�8'�#���ձ7�w��?g=b:�eY���*#Q��#�.���v�8t+p�MCi�WЩ$��F�v��e�a2�o���V0F4Jx����ajx!{�'hf��4��C�#���۩�~��;N�t��� ��ͥ�*����Ɉ}��|u;�T[�E&�il1��w�������{�����`/=#�kYKs�#&xW�j���ty٫68�������@��P�%8t��2Rl<��-1�>H�V�N���@�׬�l�[�L3\2)㬂�'<p�;8�-�o4I,p��q�2����-��}�<}Ƕ[��KY�:�ޱUŗl_ؽ�Z�2���ܑ'��$�e%���t��¿�<BE�j/��xH-uO]<<�����O���`�J%Tk�xILd���to|Oi')_ �DPtEj���{�J�_{�)�y�:D�!�>t�R��l�L�A��(
�W\�;���_��`<xD0``���}Ŧ��^G��7L��F�υ�)�H��{c���������&Fsdx���X..�Y�s=��ۤ���6\8�`�t�ncI��aL�XE2�0�9���ʚ�ci�1_-YH,/5ßq��
4oA\t
'ѕk7e��]-�� ���r7�ݴ/�Te����0�pրR���a[8���!w���H˲�k�