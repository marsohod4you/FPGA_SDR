��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su��q��h,�y�df%_�_��Vi��jP�"�9$��$F6��� ��
�����_�p��Y�M�Ow�Td�X�C[{v�L��kδy)c���{WQ脆�M�X)��{b>�Y��V�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P����0��ܴ�t񢞦�Z)�7�{���O���Y d�7�.��I��8���c���׼��U��VѲY��=K ��#~q����4����Ĉj,)l,��ۅ03���c'b��#I�Q�K4��KB. ����u%�7�}�eTB ^�����������W�|�1c�*�K�������ӧ
,�pA�v�h�K���������`%�=�x14��]�g�7�*�ִ�?-�.P���~hu�&�X�����vd��7 i,��GE�m� 4�r.�;|-�w�>�R>�dU\��2�*��֒��
ʕf~����4U�^�o&{�.�(sAd�0�ٔXQڙ�8��
3=�U5��cӨ%�OE�Q[$W��������ؓ�$�$·�����>�uQ� `�F��d�����ٹ_�ʅ�е���P�d~��@��z�kR�CH8��yk����\S�C��j;P�����S�����؜��^_��8�L��c>?�<Z�����)�|K���G�H#�s�`k��e��N�9��}��$�66["{�).�y�]j2���6S���h�s}�`,�����A�*��S���R�-B�Lն�����X���	���FQ
T�*I%ѡ����i���5.v��Qݔ��!��=��eK��[�/�0?�.+l�;�Y�%�s��p��G1�|p��_��e��u����^ѽ �V�M?#1K���O��bA�s@�v����\�1�T�		[Լ�`A���O�ykd�$s�/�@��Q^}p��qV^�F��ex)��4 +��삱8�q1���)�$���x�Mw��T)�J���c����3U�(tn�U���k@A'`T��hs3��r�����"H�
�H�Ȕ�'�Fk���TEޙ�J�h_���^d�sa�~�������Mm8HM��z?����u4��2n�7�j�R�*�QG�U�?�)$�׊�W	�9��<��p�X[���Ӟ�_��Ӳ�|}OP�o��ߜ��dNb�雭r�<����z�ל�j9��Y��Sm�NW	���K��.�� �I�!c׾�xm��bĵE)�9#�KM%�����x���qS/$�Y�\d!H�E��@�J?ܲN��ޗ���Hxv�8��M�h��#~�Xk� DU1TDN�v�0K�<?�^ǎzԯ�5	���D#�_#��{r�	���|�1:��쎙\��h��$:���}r0�M�&8��f�� n�H����7%���ͭy�R�
��oX.��4=��T�#� ^�l4���T��;�zt�¢4<���GϨ��YQt�849��ZQ�Xs�ge��h�L��q]/fr�8l��
��D�T&ȧ��9�]�q��J�~]��4'2���0�ڸ��\K%vƫ^c��_���¾{�D3��cʩd��3i�ٕ�rzG�[����;+,�9HU���!��,6FG���U3�����2��t��zy�K��@�����,�B��2�F��\b�TsG���gu���3a�SF}06�ؔ	;��ړ@�+av����+r��h��XȜi�Ȏ�)i�s�BmrB�n�'W�p�}"��uZ���<Bp��D�� ��P��V'�0���
�b�f���&�����,V��ʶ�i��Lw܋ �OOW�bE�*������
c�"k`�Ȇ�ht4����kLa�p�-�������	9���U�fS'��	��_���f�$54�0�<�-EM�Z���;�Y��j���&ÉX@�UM�"������$��}�� ��8���T����g7�'b���(��Q^לVO��]�At:7���țm���G8F�ã�9����HP_$r��S+�&�ms���`޵Z��&|��Qɭm��\�\#ݗ@Mį/y����\���|�d�/gipc�<3W0lih�`b ��M���U�C㳆ݡ��	�3��>�/?Y�Q6t4PsBz�M��O\��{�����i%��O�U�����G� ��I��t��$��0���&��1���Wi��.�P��$��z+y�Y~k�oLy��ʚU	�m�!��vb�"5�d?��5�
��#�<������� �s9�x4 ǐ}st��.�@��m��3!ue�s@��v�|���z0Io�O���-���h�)��u���Ճ<p�5Yx��A�|���x��Wa�s��NT�o�F��5A�#�_y�U�>�n�Ɗ�·�r��3-��ȹ�=#�G������hV��3�Tk��i��w+�	A�F&�����jg�}.G�I�S���aD��Ê��\�o$��^�~>��1�֙+��P�7�
e�,t*�zL74�JcPO��k���x�Jp۳jo:���]��kx�&N]W�zj2Γ��Nf<����|f{��C��M���X���厑���N��S7��e�6Ⴭ�
N�)��ӛ��t�_�t�&ƣ��\�0,������&=�Px58�F�<#O��eX��&U�����?}������ �Nc� L$��;'��.(�NS���AMP�$y��9"����9�Ѣ�}x١K���G�I�(_&�H�O_z| ���a�}���b]
]Q��;>�8'���2t>�t��x����k�T���\�	�����<%ұeBW�E
�f���|YqoN�Nq`h�YT�W˪���+EZ�j���&��?��6c��\X_m�ǣGs��Ї�Z.f��X��
���P���Z��*|#MFk�j����e2[VG0���yƫ�c��ΗE�g&�ѻ�����tJW��k��N��
(j<��d̮�||��9X���X�c/��gmm�5�T:1-���n�1�C���e���㥳��M~y�+�>�y�`NE�A��92���%9���Hȹ�^/.3��KH{�N�m*�(�؀�Q���XPP"�,^���ܷ�`@K[%�������i�H/��+����z�U�SY��^z�.�pS8����n��`IsH��L_B�P�d��{���$A�S~�iCu�R�S�����]�ޏI�S.T���g����&ǿ��֋_ֹ�5B���m�G���X�
!����E�.�������y�axn�)��1�f�H��*�'FiUZ?4�+�����t,a��f�#6��p䅜)P~`v:�ɕ|W��/ą���⁏�^�TÐ���A�,��� ������P�K�L��9F�t%y7�p�!�ev µI�Y�]�2��SТ.�%�z��
Vǋ�������r�%�#�A#�R�k��G�I�T��3@kfA�|ǫ����(6�.(k�WL�\P�K����J]3C,l��h����jIĊ�~79f�[M	�Nx���-@C�4���+^4���=�!����`"͢���_%w�6{�JI:�ȕW��i�
}/HP �������yRC^�:t���ra��zଐЗP'�^��L��q���5���:�ls�{W�����O#,��K��ܰk���M
�ƛr�� ��@���1�Ө/��RK���[�
lNEF��9\TZ��a磌-He��*p
8��Togӥ�{���U�0}R�@6φk��#���Y|Z�͡q9��{�3�z`�QvSИ�����q<��~ �F"B&��B{��Ajp�����*������>Fő	FL%�S�׷ _�|����ܫz���À@��a��TO�ލ����<��ŷ�O4��k9E�@?��Ӳ�,���=h|�BR����չ0+�Z�v�*
�}�.�;���k%��;�'j S1iGk6y;?z瘭�ZU��C���7�[�1�H�.���S� W���舲JhI�:��]T�Wҫ Ī�:<R�mLO��0H0/[f�/W��� �����F�!�aӝl��&�X�6\��5����6�c��Z Ckƀ��㩽���C�Bo��e�30�p6ַ��KunV��a�A�%[�l�5s
+U7LB`�<��^7�/a����9��wܷ���[��܂�$<�v����Ât����`^7 j%�U<Z���B�P�z��n'eo�<KHf�+2�`��N�:X��=�?hluތ�;��c���I�����~:�蜭<:��R����1S�a��k#�t�|�`wmj��)���VF���g\e�Þ͔.�_ �L�_~��X}O�:�'jT�?G/���f�N\�O�p��(ӵ%q_��p����� ·:Ƈ�-���Z���!�������%�&+ �>~JGv���on�~`��	9�4pR�??vN�<�\�N�N1�k���{Y?(z�)��t�3��_{�r��Hϗ\�t�d��@�T_ň��F�s�r_�V��u ��G�4�s�����C������[���z�\�	f֢&�i�X.��^���� :,�D˕T톕9�5�@�{��kj�Ha	AZ+	:����֕�~^��{1̺`�9T�	��:����̮�9te YM��<գ����eh�^��"O������Rd���C�X��jy]6�e�v��!�
� ��$�7�n�bc1�-����ŭ����Xȍz��+L�=�)��j;�*��OI��;0��ڵ5��[����h���_�^��dѶ�@p�֑��&��C�-Im4��8���AA��9������=Ro_��{�	� �sIV!Y.m��Z2��H�9e��FaнL�D:�dB!�R�J]���ؼ�@<�c6rh\Ǣ�r���.�7L%2�Bn����]�J작�%��P��D��4���� �׉���C�#t�*�g����X=6Y԰[s�Z
����u���J�ai,̜�6P>Af�ԊU����{�ƶ���k7��)�[�4&��*��4��o��&���ORtMo!��߄��댃-T�[��į
ΤW䎥�c* {��h4������si��n��S��B8b	;3��"���-�U�����c�Uh�g [�Q�7t�T����":$ȋ�'���7d�+ Ṅ��,�U�e�C��6Q/��c� S�λ�r^�����^X��!�n)I9U0���Bp�D<�yk��E����!���YB<Qo4���l��,˴�6����i4�w'΁쫬V���< ��I�Z�<��}��C��M��+�����H�R��}�>9���/�XTs=z����܎m�/�5����p�T�~9�-�3:�\���-�����Ra|B�%X�~�L�ug�$w�7r�3fM����2�E����ה��K�~�T�v���pZQ��y�C�ͫX��mn:�*>������'0es~R������@��u)�n���d�H���b��i�x� YgK1��h6��[  S矯�XǺ,�L��fO��0ƒl�T�����qm2e_��+#������UX����3ʮ�F,����[�Ҿ�����0�,+yHAx2	�׵����8]��wb�.����!��@U��x�"t��LFYÃ�#N�8٫�������6=��q��~b����o�e4&���c������C�z4 Is�������E?]���^3(~����f�ii�;V$�2=T�}h]G����yIS싣 ����~���3��=>�ь��%��J��)���j���a�~t��{E�"-�q9�.�\8q�ĝqP�I4�o�%��A��+N�1_,�7�U��2=���!���6�)8b�=���đ�h�����Ĵ��4"�F���]����H��	�/��{X"m�H�[Lܱd~�Sif�~�;
��l�4��J��wtΔ'e	���[�ӌ�-�NY�fyO��1�tS1 J��}j��qj�� �E.�~a=t����2��v�ɘ��������>Ohl��������F&ޯu�r�ַ�*)Q]�r�ٛM�a_��F��M��z���j��"�&��jJ�d-�M��ڒa����%0��-��Rx��-���զ���3�R-^O��F#��V�=�:���r.�Q����,o�{��Q��#6 >||��꤆��يS �Ȓ�6�9�b�DT����� `�{����X^s�dN{]�1�j�2#R�)�'DbRCSS)|�!��+@OxNmfPR��iD�TQ�FJm��j�p��e�
���2$Z#~�\���-��^�������t�0	�׽P�%����M�o8t
��j�3+��JUe.	E�%_��������s*�7�o�P����ja$�ߒr�%A=��B
�K����ѱ����.R�dDK&���.v��k��pj��������<��ȯ�)��zU����Ĳ_)�tHFa~����__��m��/I�$Q��(췤���m��2��0��
�CV,���!�ᝇ�6�^��[�J&����*f�D�J�t���P=9��